--
--Written by GowinSynthesis
--Product Version "GowinSynthesis V1.9.8.07 Education"
--Thu Sep 08 16:32:32 2022

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.8.07_Education/IDE/ipcore/DVI_TX/data/dvi_tx_top.v"
--file1 "\C:/Gowin/Gowin_V1.9.8.07_Education/IDE/ipcore/DVI_TX/data/rgb2dvi.vp"
`protect begin_protected
`protect version="2.1"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`protect key_block
HEBaR9vWIx4Eo9quu/NLtUzICJCcQG2i+8yuEC+vFEfWe5r4auq3l/eBJeo4ZGdssj/RX6qzgPq9
mrq5mbA21FfMMFRcjbvFoH0VziSZp0Zev72JlkzGtsQoXf5WfTvqAoOsqgR2dil9OQdtpPU9P/3L
Vfn3nIXBTzRXy4LcTwqoFDQ0V5HyEmeduQ8x5VjiD+V8dzCxIGIPxOpwSt2//KaGGyWDYnxuvu/Q
Zs2yFPSvIJyo/86qeUwiWhZvca9TUbfcysaeLL2EmR4yrsUAJ3aiwkY567/AMsgf59lQC4zYjKLc
7NmxeJHaRZ7QnIF7r8AgqYYdaklwD11nuzD+WQ==

`protect encoding=(enctype="base64", line_length=76, bytes=67248)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
pymUK8zoCvcl6R+ogNSzM5MeeAOrfOp2k2kRjVLxFrO4W0HDzj1DFDJGUOGKkfhNM6KL6J7NNSUj
lwo0NIlnt8SLkBtgep6D1DYPwtjrhikMQO0UGVT0PZEpW7Psvph6zZKA34Xy7BRH5RJ47kXjpi8X
Wz0PVgJkveRswInBMcNVC/XVhYQpRS2TInDqHUJbXyNTIlPmtp9MnEuEqNqQPn53yro20DCPakBo
xHDEdoBtTt7UWc91pm2ZLEJTLmJranjsK4p4C6zKyVACyrh+sa3yVrxVqzZMtDlolZ562CBDNTU0
Fw4eOCyaLMb8rz8dbU0JyGpGVlpk+4u6pi2FkssMFT54DRn/7NJm8KSmYkVpq38zi+2OfBbELXCA
WvLNeilOKYR1rXz2QNxD+ttopwtceL1FI9E+/PQoi4IcShaCQZWJPMYiOR3DVHM7JlRlLeW11nNh
PKgphq6AxdW/RH7d8qYLrKbSnmsJFi2GqZbb3zkeUpfpo5VxZzXeCYfsmrln+4RS2DtiITOuNkAC
P26fjgR/mMUG5UJPjzGg/sZYF/1sWBPGvuqRKIcBf/doQYWxkpMY7IIuQrxNZG/qUqNFyqVtWsti
4twy4SKzSzxXV6R+WOeZQNBVojG5jUL0ryZIOQqXzcbfBeKBE8Q0lJo8qFKPkBhxK5t4gaZSBv5F
qHCTasmHypFMBMxbp5gT03npGB5uL1E5H1gXjYu1FjZ82YHBvfx6vG1Ny1Ca/l3gdEx60mjhGsBY
hpKfGTxy9pVtQpTDr2+KRCPbGmE0k+ThDBTrH6bLxU8v/bLnO1x1bM7Ph9kYcKPit13UtkphAbBA
JYuOu7Lh/uf4InZnk+J59YOIGXxKXu1EOSL3ws6Q7ly0oOTms7qReV/Bj1zqKpGBqnXS7fcJyJrO
M4R3qhhLpBis1QXalGcuotXO+nlU3SMzM68xlaTorjpnOvYYrvQ5bUQjCj/L/P6cmUj+MLz7djoW
YmjRY+kZjO3JNOq1XNJimAVYpMpRafQpK6exLxnfbAmmQmQXCmXU0+sjC4WF6lNaylkcHqO4rCfC
XAz0l8IjFe3HykGGnqElRCb68aEfQIYt24YzaL8p3zcT1a7oPjYyY9dwCE6HyVrfiuqUxwcjUs2m
mbJrLCfnq3YES7ceCRpudC1bjpbVCiBSIntql77kzrbsj1la4Fo0wnpbcQlqt1GQTTAPhpsEKYd9
iXu+CQDx4fuLbqBq/fLVbyNqPMS0tFL3lPecVO6F0z+RC5ZIdbQONKuvspUiJnYUrzps8+VGsM7I
Tjb3laexpnjR4j3n4Yu4HVscTdffhyCcv2jXgT3udYlpCKGtUd6GI/aGgE2nwys+LnBOOgADofNb
HKjCsaNKu4D2yUAGI9IDovdGqk0GK4d0XHBPrnh2qmYN9AjZ8tfIOl0Zz6z4g3sOl0xYdPnkCIl1
zLQoh83l9lX8PG3xTCDrt1OvPqJ/Gq6Wt6UcK2Z6MRXZa0B/uuFd+b/+wGu/v9etNPfrAASRBPPH
9T5tSQ03UR8FqAuVk4rZ9BuurbFhP9mFS5FY6knY4iLBicj6JGRdnIw3m3dDD55Ky5OqBhhoote0
obOxPfKpfOJIi3TBE3hTWJm38A8yFJpQ6tVTt7ksQwd8DUdyRoH7XVc7JJaIBqZKQmtNLp3LY3nh
1XgBikD6gCScwVNqpF2UQQY0hS9kSYq95r+DGtuEuWHBk0s4kwyo5iWNdP48pjRjIDC61FfE8bLS
9o3jAJ05E76k4B0ig3VLb2gnD/6+BSY11FaoSKartAfHy+AuTy0L1XAVoCodmcRcrbAibbhWSCHj
TV9VlcNga6BIyiaKdBsH6OzXz//B0X9jEiZiPdZxUGSFbOm0EqSMgMwZWFszFTp9WxCRcsK5a7fs
wd1U3JJQKVyM+5WoFxvujDmpq8gx/nKXHHQl1RJoQymWxUJM0bc8FK2MO1wjZk5+mik2+nYVKewV
/NOBtw6gJOGi0tKreC6dFtizVG1yh5wx5x0wSPcumy9FFVdkwLUyxHh1kEaphwB2L8S3LBknRV3N
yJVxHPnhioPhy+ujhwqVx/9ydVKQMNAO/6p8+lYFTHoQ6tVHXQW2DAVyahBaMZDvo4mBe8vSjrjJ
vy01EIB/xW+pDy31GhcZy0dSIO38MV3+0/hTt2HKXV/jvoDiE3ThFFfD9smBFf7osGenuJp/7j2/
6eGOnZiLTGp2XxhRLQMeZYtAVK3Q2liYwDbotfToH4Dr4dL+2JukypDjH+Gj2kL1CmLJ2AIOy8hj
t6MhT1sWSdfYcSMCI6LBXMQd8C2HojaOYGkm2LlBaL3kq6XMKkte+noArifV8AYuDLM4bhDowIvd
pv3CPmtCgiMA1o+BhvH3WjbMejeY/kfPrRCGjGRM1A9BYikuHZCaAv9OyNMw+f1qU8nMNYBvFM1u
IhycPEfg3xbkptmAre0w7e86yiZbrCpRuC5tDHbkR/qEfLyXc/6ySbhuiHNkircQetRagu8bC/Ga
9aD7VSdTHY3ViJikIRnF7zrShb8L2bTM6DtlDV3kooeDT13tycLaL8KuhuIp+UmX/da2TfduKQy1
kCNRDeV6vEAlhT9EFZF5ywrZ5GyNAauo1JUt8nUS2/IRT1pP3eXMso471/55pgqHAdKXov6a86FC
3YV5wbukmHI5PVzFNZSe61Qrhh82HfIxoWX7Cj6VrEoegBDmUfaJmYQ54Uqkvz0tKwPBj7osXVEW
wzuUAW7q8K6XMuEQ60EA5TXngF1aWPJv71wIHlhtdaSuOheCYLCaefzRD64rvcdjrIGVBtgpWCAA
ukqwomGkH074umIkcNpoO1EGAp7DHr68kiqlXbCkqQo//aEB5t85k3FmH3/5sajfxmfa7VfrNWQO
H+XOVy189E7EopDadtzP/QSWAA50TTVWYSizp0MYlMEeni+dFM6+ItV+rn5l6Hr+BlDhFZf+/GaA
yaMeiCvP/D/9SFs4qI1Jeih13/VA6BvIi30FyxNJZza0R0lDgWU96q0QdIOXZtmCOfizzSLBTTbX
dTVeXNF5Ky6i+/iNiTdBx1Vg4yYqyENqQu5+i4TifeSg0ybhihxjG2BoKga7R5MGe1ej6dAV7KQ1
UfiNVg4li/Qk7QEN8Qb6guL0oVm4bJwPRkHCryFPalRTNmUqNMKLKGRrZ1P4Bw7+GpdWByXGbmJb
+Gyvu9X0guKB3/DfmubivcsjVoJdjhJnzj1YE1Qv/6qoULg6evAAGvlwq+7jMngxYa/aTrb/9332
jSxofOnjxvvQqYOeUR8tTnSeveXvmgWiPYQfJ6zCM1fH/26xJjaODkSDqS2xdDFwddVjqEZ4othJ
D8ynkG/CzAVbIYula9mCJv5kFFEVgmWAtBv+u6T9qC3KKOTQoCRD2yy/v8rHv4TFSqQIbW0ybqxi
goyVw2tqG7d8GGkqdshX/PIsWDiY588H122YeyiC7Q2uHIPwwz3QxEHV17UbHmAdOzg+9Cxt58EY
Lq+XtO6zr9pM45LsYuduRmj+poXWrxpN9icxfrJSRCLHEVks2mAEDd/lLinqYbJzyx+d0L6f1Suw
PLt9NAeS+L83G9shCACJqA0izshrA/w7jX3+kMJZ8W45jG29dUnxxqCU6oUj1XjFb0kCY1/QRGYk
rPELY41pUsxX5d0Ak47a/USMKgVxLiwNtiWdzxNioYRepLcVa489VaK0A7GQLGNBCm0RTOujhZ+6
dc4zSXS4YsI9sxhTwrrieXHRZjn3baYzWD2+D3/D7shYDvSlXp/xnN3xMvVGQBF1qUN1JgrOGsSs
nuYnMjeJ0le1cUxiYl8QfaBeJ0/X0N+LS84SN3wfrDZgMV574KZrm4AKhdKcGR8YtV+mmfjRgKFh
aNYjT1yFGG4I7RyoTvX8HvWEDQ3GfDj0rda/qbBLdRFcK3SPnTStDR2fBmj6hOQ+jozpxUsEdB+k
33eZ+qvPNntb4BoHPYxJk4f3ay9Xte9lupm/OKtNNj69oPYuMbaPD6zzGR9l8wxJelBEXkmMQVGn
iIjrX7R9/OdzPoW9spxChxRT7n82fraaUaHrTbEVCDNaFq/7L0bL7CR5OmVPFCcK/F4R46PxvpgN
a6+pkqlUkrUuSQxRqa2nVUvqRne46VhX6Etdx/e3RTUGlk3hPuttqkMlLLLbYovhfTLCXPlnaU2U
nTkbxLX4NJdQlb6oZfYaTI6if1/IlnVcqqkgbteDg62SfpcPLwsUrDlIwGRUoainW7JZyAITgs7m
CQ4EZVtH2RzIQuxahsEbgZGJP0yVXk6RGgrWehel5rUfI6Zt5Y/ly2n8BrNoPUDUplUV9ifZNbLu
kBrbLFc/CA24ZBGiDKcYDgaeeErPYEdcnczWqy9tgEu+rZmGj2e28Lt2xHW9xjs7soGbqlcFZ+Uz
Fb+YG1+1aTSqw3NU5vUfx4Ipq/H4rFaNribyQTsM2e3SOAAeCJlM/cAJQYVGZhh4d/jXHA0J4Npx
izmAEqFRaLvEEYALO7V9RBKxufz/7QDZrWFqpSSeItROmcfOS6TSHl0IAZlOGW1A8Zh06Hp4G2k2
hU2bdOlCX4OO3x8t1DGMbwWfZX0JZgmsajRCXvOs/iw6dS5dx6Y0qUgsrYNu+6Ei8oaTddiNqyeS
Sx1m7CPO6yrNtSh+gwwfRE5Pw/LVGiGB5J9ehSETXKVlPyDgi+L3zKSe7OWH/XWDRzY1zqjYW8qg
rFLauv+ASf2W9rnBm3xBSV2uQNN6m2spAgGRW3jfw8lTV9wd1/0Pq/yAhRdFD9wxv9sExXbbY4vC
NsyH5iK01Qd4w6ozLSKp5G+yJhNdVQCkjc3kwuun7yFSK9VnNcIdsG992iWRHp94Q8vi5MA4EEXR
XDssdwJ20meeAxHl7S2D4fyVjnvM6kYN+23CZImrssdrXk/KO6Xm4q3tbDcgIyVzUmNnyZA2yWVV
4lr6vHcMi2LFyVXD55hXq+S0uegk3AIdYflI0K0jQ9g46ysbnIwxeDOCz/fc45uTcO7bbXwI16HC
PSDxPSjjVaMOzPucwzBa9CCOWt9eXJnqnkMvrW5oYmLGIMaI4L3Er3sw6oayZSmLKAfqIifUW23g
fh50/6lESBD1aTlpZSFT1getkxHMb/ie2G4URuxwY6q8PtAd9HMvPcnAnzjGa8IcqLqSY0cMZyvN
ggS35inU5GkyCuz1bXhHYLnZDe/XuscDy7iD/cFJmY9cbQbtAi5eS8b7RoFRf+QY1SPwOyPY+SGY
pBxz/YHwa9DkkXJRTTY0NRrrRq48o4jRUeSfiowDEB/upN28gN2iq6iRFcN4rvWM81W2v0JE01r2
cP+Nr0SsBSEvnQnenj/cMzU9iOodqdJsGvftiPAmZNcLmFmEH5htbIAxF5vSymspd5AvT5bUYuKJ
l4M99LtrYz3HYQiy6SdyfAuSXVCxc5Lz4EQnXJmvudnwIMGXEAUaTUbNiKqv2aiYwjoxR4hKTZD3
DHgSlZCs37eVUa0RRoLLvujsJ1el2PuKtbIHgzicOQunoHVlOdGvz5KbxxV7daB8BV+DlPPg9Kld
E7weXcaTQKRVdEN1oUWeXm/txJYV+ArGdEUA/LahLvCh6KilTH8fC+I2KoqBmucXCBc+LfaOxPXa
iv4/3hRgTVHQFpADWqEDwiCH1Vae+Am0IVeJ7U0LWm6MNe5RbFCZgB4GxLTNtcBvylgKouEPF9ol
fmnZdKFZhNk4WmrT1M1LIgtJG3Zcig4FDfE8AT8Vtcfm4nbyEm3cGTTZ8qUVBrLDUX43EnO3uRNZ
EErwfMfnf+wG4uAapPRGwLk1koI7h7R7w7qg0SM+XRkmdhVAhkifAebtMuLlyubhJGFZe6LZtpq/
pTyeQGTHrnVKX9+c4c2MMHxsO0NCaqWU8/PqzSSd8hgarN//IvlTnSSpPEMAQ6R1ikfqxr3+x0+p
ZSMli8YWo2TBVeo0YUYZ8PxYwf027Haxb6lOGz+L9v4b68/yqI/+AhAjM7ntngZyoZIMmAyyt4kv
Uxp/9sN4hbXziNbzCE6S40zaMdcNui4/c4baV7jskUhRgldVg6QG15df3d2BEIA9EUzPLC/c5yK1
m7A+oByzawKuiZqQVMDnc9sU8Ge5nX9OudSgafO3Az3PtBhXWtU548ajW8IrLpv93v45H5JBPrUh
cW44e2exvH3dITYwe0KNn99d7+AeTmRVVawjVc3FbfU3/8fthLPCPaQBCDWglqlxXUcGejZOVSZ7
H/wHSqsxyQPRuJE0tXoPYfJeW+pfRFytPx9ZNYyYl5l68w7wCWmxO65dpzHZWGIpIi61pH0+uM/B
1LepXomcXzgnwkJYSP45oPtPyNP93QmxSr66hlv+aX4RpZHzYC72aPUDCTp1BTz2drBzmgzllGDA
hDYKoZdmeW8XVdxSYnhfbCV0NSYLG8opqH4cMljvYdgMxaJ5/34oUQyJtgjH0pDNuhcz/M65Uf8N
2D3ENE1bHTADjrCJR1dSzevJbL3VOP5sU9TRXi17A0Els15NbdZo92wPRGjw+DfLkX3PJdZHPT9T
+B7kvj94/PNleRRTHDxQVxfra+ms0j1utF94foIXLCMaQ/YYuE2/OkhN4HK3/VdpJMsOeuaAOESK
ri7SQH1tPqCwlL+UyaLmLtbJ8ZrV9gpowc8AMfiW81XH1DG3Gd/NEJhAuBUhFon0wsZWLQiErR48
BkqCp1XfB4ylJGgoNooJWVc0tOQbLyOscWhbvce7o22vQigkmZQnymFgzrHE/Fmw8NHMfnMr+oO7
EQ8YLd2mtejf5G1iDaWNkDM7MB8MBGL9BoFZzQDHB37YEiuMDz/em03FhexXNj8GPUB7hMZ1cETl
bKvY4OEUDhzsKNbpIlVQngHlHkjKi6Wvtw0RFRp68q1iqmphpy1t+y0TOJ7RiyXlpE6r8mrL5A6c
aNInpjBm8L8OutyZhpsg0kTfjhu3/CXZ/ZyT3uWTUh1rjE/qxxF8wa468erlgdiHERobkDbQgAMs
nFIDTfYpgdcIpopNhJAQlVQGF7Ug48bAccCR3LO4Pr+bLLuMYkcFCpO9JHugo3neGlIgyxkVoudu
+76unlhYjduCO2SAHMh6HFoRSoV/8Rp+/zD9Ne8tR+cgLV3nzFOJENWplDFVtpWlnQpz2Q1R0GIC
KXuL7LVwg+Be3o3tBAZLH7PTfp9a68VASJ/i6JG5N5jsc6uPhuNLfXnI/MPrfP6RF7LZ/+wujhU9
RCFc+dBAYhPb0mngu3K0UDL79HuHr7+YYGqMq8zBE/xrdLVDb4u/rN2Ld9cmVbcp+3YDNQRkvrIn
+kI1nCfr7L2IpaU63oWveHyl8/wORXB+6VzTlOFPfkJ+wjpP4h/hsR9A2qoDahV8eXEbgh5PWBiE
/5GCT9lz4LuqGBUuC2duHUa7YoOWSX3JmvkgWQ6B03AUHma9RO2NalM8bjmPdpPlT4TBkQmm/kUK
rud2zplNxn9+dGB/dLi76TERba4Y8HjBI034PYdDEmPhEaT05Xoi2cS0yB2Jz+vx4Qi114m69yOH
464EpI8oAr3HZKif8TK2pswGyzpFX6MQwCZ/kEau0JcyFk8nY+D3UfZBwKgIDtqoUZnLSKFgZjZ7
HI7izgF0Otgt1kO3ku5+r1NLbPjfxgwTSHd+i/wKydMsp6eSDn4yBPBt+FIr4ZmwdJNjwh7HL0Lw
cOBq0hOF0+F3lPGl14KAxW7BWlKaDq/HjAZz+2EnlsxxL+o5TaJJfb5QXjEExsqD+xec5w+bNy54
K7Br1N32mMmoPnd2DRwwrhfyCCKRoijuNBaUELBKdFOMB8unR4AV2WCJen3XOIuUyaAX0KDl4K1W
y33wTiPb7Qcjzi1+GiWD+ppvVc31+IfXynKG77cF6dOA6lxwxmdIlNVEWDDpElCMV0Zry6Am8t5K
UXfvHuRjp7kEd27oWmN3Ged1RTfvEI1sy55ZjdKVqr+StnN6cj6G5ciCAztLUikV9MGioHQqlNVn
yNcorOtyqkmPyJZKUqhT18eWrUAvKsHuyz6jtnmzZkW15sjZRoWzBPzxpDWxwCI/uq2AxJF0nxXN
a0pbFGu3+7jV6m1sTXWmS7fuBRgtGeShRkHR6VEol6l0+CIj0L4fBNrRZe4aSsnpKoXTMUwngWFC
OOIyEyDR1urV1Jr6KY39LwYJoKlm/TvzcO8jLDnohzLYiFxJ5uKQOb/zlWrScW9/ec9v1YUrlI43
vbhjwVwjOFbfu61+llepP9JgyOZKSQM5L+npLtdo4BEm+pmBthdZFfImBzVxOAyH5T6ZlQOTgueJ
rmQTs35JIQS+ztB+nJyVrhDm9ehH7+CQtFsilv9czW1jDetDY6R2Ksj3j4CK5KFw2m+ETIvZSnvq
Lu5wUM7kPjaT2FzKnRRLZfdx9nkbUK+52FEgU8SZppBt4fpsMfYAnuat/IJqGAw7uMJX5Tg/oOty
3xqvSb9za1jvPh13QW8lN2YPovq4DLs7vq8FW90KoyZP7KmTi4U9UCHno+PUauSnQfDrhfFaA9Yl
rUu4bE8hLNqSWibBgDfwc0pYT2UTzey+vWoD3UAzhbsx2fP4gvWnvFagRyi4bA+SIsmLdRo5uFQ/
/7TjLXyeCyYp04WyTBL9WF05+IXezn65GyXGR9AF0EcDhjPPuxGTe3EwZ+6oeKbnqH2LZFAfPjew
YDNHJyj23lyojNA/y69Y5LsihRK4Bn1jWplJ4EUZEruJFhAwRf2l+XXJg0EtvoQk+ZPlortQ2+nv
04N1+7PSrLMeQaqTgn9Xd7rkwTTooqbsdH3HJ5p/qerAMxVY1SDBMZH2bprwZ7XP2QlxOa8WbDJv
gdb0FiJABI7JoVrhbHwuyc3wCIhu34xasF6xPZL8tz2yk+C4zn0am4/nrWQr9DiXqlPoiNhP+EQX
MKsvBxROYKItksWCm8bpbEATTUlX14DFig9er+OvDYMl3vQ2HYEA+hKHfWtYtXTxG8pHRGCYgW4H
KwYExOgATepeOiBDaI+a7EVYTBrVqKorlClFHUumnaQMAAdXaxDAiWw7sz6EBK012A9hABGdD5Zk
3PaXV++2H/+tTCTJJ5dSIuQHavENvFXPB17DiO58LlpaB+CxAix3DBPLZXXNaWnh/Md2QURp6DdW
b/slsC6qze2MSZu5fgnASHTXIwmhh1vzucssKQBaDhr9Ok8NrtC+UKHEgLr2obXnwoL9ZqOc388A
Iq7XTeIjJpVTBgeyZuBjSzYpGoQUZhpK/LMqSvReaAaupQ/sZ7Uci5ceuvBArEfImwgmPodFWGCn
JGwMn8P2+55IEpeBqOXc1Eo3xkA8yNfY8p9WHDu5MHeKMt6YZI7yUxkfzuFpC31MZJUr9UnisvTI
uPRbo0POfrR2Ax0tjEYrKFuJRXQna8V5bxHmEKu5c0oty00Amlmyi8Cr9f7EzvtHfKH/RAF7t6xr
V6BjwzQ4JYsgoM139UgonaxAhswTl2PKMY5fQaeR/hm2CwTDDpVjVb9u6MKEzzV9qSUX0FUSZKdn
1LmjI7naSUxizc4+8eQUFtLuQ2LNAGeh4jkZ/qW6Lc3TY5scoaHfanyyakKartDLc2Sff76HnkIs
WnQDp4e2Lfv3j1HRlE/iASgAALpOmRKf+7dS7aE2EqN7auW+9EpsFXw9Fs5YcZQVEc3k8aD8Ng3A
XrwBvH2oKvcODYNdy1F1rgGuJjfd1P6d7LLE5SSGvNiQl0u/bKVhameoPZDg+Y9CFlWaRt3G8hpt
apIcL5ZR0SZsqtDZT7BTGjZYmVTbR3x5nkMZe7RYsY4VGnGeYeusA2f8KiHRJ3l1pJwoYgwRT6AJ
QGaeR3OaGGFjWZunH7GvMayg4cQ7Tm+dcWHlUJJ3eD/5Dh05lDJFN/8HDFSyUpl1pU1yRyZF1e2s
SA1m06XX/SjyvuCinYDOUBYLTiQtJ+WyABpwXIBNUXwu9U9FXTdYJEQPGJxR1RYWP9FjlQgf8q9W
hPQ3J/Me8TXZiyhRPLPGHuWN6GknNrNIZy9hK3ig7cGhYjzlHW/xvaHn3h1/5fCohe2uwlYAbzxJ
h6XgrjHAxxG2O/S+HXCudQWRhkmrXrN0JME588wuVqIy5dG6+eLp4ThX94gv8fgGb8KZuE71I4Bp
nCwk3M9oE4+L90c91kZa5OIEzM4S1bzsI7/f+2Q4LFsbrK0CI3MorTiIFrTJRrfhlvi9lMpsQ4Oo
ZmpIAy+8RSlPXhbMW9x3o3FenwuzKRIcefOIuywA2fbl3PHmzO1oUpRy1NsrRXKF6R8EzaJr0uhp
49GgrYIpKeFVfXDyK53ekxhjJp+PuaP2FdMmHevXJyYQoC44ihvqcPUkgA7pRkT9z7CNZyPikr2K
heZMQwpmk0vz9aUmEPJapQkuEIMkSxYMPGj8nNV4Rv5bJTwXorYM5c2jWeBcmmG16T2IN/Oa50Lo
PxpXL+SQBBurxFAxNjY1N0nv7NK23BhGBhx+9uKNM/Cf+VTStDXXMTCrnwSoVEB7M/to5qdJzCSI
7TZwNuag6V/WLulHzRejfeU7/9mVl7NX/rYd9NdxhpHRJqxp/iaw0WqxBWyl1wUUjpQATmSCkT6F
cu7eBNoM4XwTdYW/nJh2Btce8WISsaNH7T7GjbIUQcuu8ZqXxB4P0ObFP2TmGCKqHaBmNCU9m6zQ
w6n1Mak4gP/WOylccEzLQ88MVSUC+Eew8bITKuv1cu3XEvsAHibW7G2wI58hprqRshLFR4u7+RM8
qb8K1tuZiKvTV679XVDmQJxfJHkwk4QCxIBtJfCCo/gvOGVoUVQ2joGvrvs3Uk9XEQBAnGg1VdCT
Qn3cgB8ueLF4zpnVe4PHXlOLnB+H31daxxM/0NmEKmJi6pf0hgYuu7lywXHryltuB8GkU58X4dze
Bl9P2y3iifygMAM2e1KRHoklYM6tr74izjSCLjhHs2hDYqst3uakCPQ6Tmn/p7ZoMmtbM9jjcAQq
TyajQPk6ws0E6gSNQEF/tR9Yvuh0PVf37i8Thr57djfVAeJ5OGvxSier6zKaS4oEOwVx7uLUeCHS
5ktKVFup3mvrrlZW1pzzSfLQmjcVfBtI0GfiXSMSvTVdLUhDRq6xQ3/j7zoo9P+X30fR61m16Gnx
QDLDmOp5PpShj5jKKtM8LFAD8xH/Z6t7zrVdYW0Nj10N1FtJOvMycvbQ4n5eY8oNkiwkKOnOsL3E
Ms+vHH/AEZrqGdMIGyiZzXK6jQ8+r1ukD6USYWuo9H+qbyPgHmddeQ2YzoqzddnIjeySMJNU2bhv
CzV2ZuD0Py2Ha5rjqwkXMvHwTVB3RZxYCU5fgsgf0OAZvuZ/hD8hDAuc/+s+5QGRAKp+6axpQklq
/i3eMkR+d21rNtJkSNxnbnk6MU9Lt0y1U5aylJniqqxXOwdle4bdj01Nf536A7WP5M0fflH0AxnU
oRQsvD8O7yYdAhclJ00li/djkbpJ2Rhv5N+8go3EFSRB9adgJugqztVpKonu5Iolq9D2cFYRr2yP
ViS3Pc44WbAAKpp3X6K5ySxlzL8skpvJgzVz/1kTm15mI0Q5Tv5sUH/fF/oLCuTJplDWM7ut6Lq/
2ZwJrGVcEk5PlrnJaFempcFzXxPKrfZRO5JK1Guczpq3I82qcLFuV56ehgm4KpdJLdCXR7O2clqT
+CPtu5XRpoKLV3w9fMsn3ciAuj5EStQc8Xj9g2FzfdQxODG39h4GNqPNf3TZUtUACmEVfvyPxxT3
4vKhcCIcz4Ls+jigTmewVLOS5iqP14ModzhclrY6PiV9fh6qYEAisJow/EJ4N6C7K3qV2liNvPzi
xsnv/NGYbJHlYci4ggyuQBGNu8LRgUPxKB1yxtvkT0d7aX0AXHMF5pUd98UNG8kGx+dkWv/Y/bTn
OOiA6UivMO29OSKOm6fOlmI1sGBM5nwhKyYgGWBKHfbn+1fx37iMHeSDND6fPj2nUDRXtkydWkFl
jD5eaAqgZLQ0H/UQ6hlpwOGerHxYf0GMXiNnOcvn68+VNil7Aer+Vdt4GRgNAEzoNtHB3hxLSu9P
EsB0efchOFGUL++QLmSkNQ/Xx47jMppOUncsxgt5WOBLwpsvHxeKPluvkliJnFuszzg7lVLUS8hV
m5yyUYwHD2pIyU0YGsuMWHTRTIxPcYxNTzM9jH5FFJBF86bFWtQ5XIJpfIEucE36yfdep6P0r5FM
YFNVRVZDehgQxL3a6zI/ZmQL5OVUqs4QNKPCnGrCHWRu4gWp+ukj0bgeFDnwTv0/fjwx7/mIS8m4
3yXsYGZrbuFgnNWB15+alVb0gpym89OfWZJ3Sp1tzyO7uYw9sEXJp+IwteOIPkvjpQio4LXjFJ9N
SSG3ExzXg6EY4dNDcrnfADNbOugpdW5EKrgqa8EZZOyYF3nYUgZ1RjZTdtS2gibPtdTAMoS3p85R
9jaNzt5DdhS2DnSxqgkSsnnce+0u0jYRsAsyv8MXrujKm1P5StEdLpOnz5sjPyqoWFca83Aze8Tv
dKnMGEIyfJ2YfshFcjmEwKV00Xfa7IUEnDtS3JGzFXOsW+DDRnQWpapH+c5flDZjXQdDLQXHOL/S
iqnqFrkqsMaPUbLRAcAxuGxGUrmhGpMNzDTptFOSYS/hNtzpvGj0f9ygnEYsowTjPgPSsgk89JVW
HIan/B0N/gOQ0f8y3pYUm/qAcuzgOcoX90ujKQGLSQ2R9WmICDl5RjevDI9EFNHZj+aMd1kHge5x
CkjC52FrtB5UTmwQda2RDYigMMlXxn4YpoikQdEdMZbj1L07DqVSXsBHt1qpnAaJlTJjUaSE7DoE
OFeN6wABqWLEG5yHrCLeo7QFPoD70WO/n9YXn7NBYRjIlQSgGr1vXZstp3ffdHEJ42bUmq7HmZv4
tz74IsomhryUU+ODmAWH+MfHGnEuAiycI9FBBVt+vC7yDPrME23jhQC2fsLs9tVwyzREtB+mQIMu
1RdOl7q0edwhT7dt+6b2r/pcFFwcOukIOcmvnSyGtQuMakfqx2ZWSxYo2ltZYgHyzAIP5lDOyySG
vvRdqTs0jKv8R2oLoIPbY2+bEuJk9C9RX1fHCcN5jWsnxPqn9PNZ3xFfjzGCnHQZP1UEP6T1BJ9u
InRQtS9IClwGXFg75EiMYmIZRHsamdauIwhKw3WAdlUGqBWZRoLP9hGHDlNyp7C7W8/6evWBaYsS
mSxp9SOBjaiViT7Pq7wz5QYcwnpNMGRjWlvLsP789OTqPT1WX26gX6WBwwZvTEfzFZO7IOo/gJ6k
llp3z5asCWEL9HCn8GJmQDvTWDZcaMwtNORf0alhEmX7eOhNujJQV57+EGjmRvy88zVgoo3try+I
kP9N/NR9IZI10UXzifYLABtj2PE7MTW/PJe+fhr59MYWk/a9IYqktXEoTtH82jC0QoOliWNtQCEu
ZuuMPsMp0Ez4HgRJL+IPv5xoBQiNqx0Kqg8UZtgSsK/+SJ9quLl/Gmv6GYsU1b8aROd9cEuHEhLi
ra+W/GyXBOYsEpXlVrbfc70cXict23uVWEGZNB0Kv3PPbnGL7LGOD1Hz5Wm0vt136Z5Qz2NqW89B
jM/QMAuG2a3OdxVjkNAlvUFsyK//mN1EPLimpbfq9LajOMK+Z3lOSf1LCpESjZHXSH5Oi08HXtN4
/Oht5PVMR0oVnPy/JyiGURPAgRulTsBNj/12BP+DQCFhDVrbhncWURlIb3dt9rfeaOtAr4VSoZ7Y
NytMfsMrU6kw6NLaDiTcEb8M+Uj46SHAgahsxA1kkYc/yb+4vXGso50AYhfrpJjV6LX1TfmPutUv
jU05vMVa6syKvORSi/jKL3gWdGQMEAztxcUyRIrtgC4Oi4y+w8+aHJRV5tvkzCHj1VYJnRK+vATl
r5YHHymoXLlIsZ8qVEPJ/JskgWywyxG2NIwv3ZxnDoXtn3UZP75jyVJy3OKl8zZgYm9nkWQWc/+K
oXmxFelVY/VS0hOJ+V9GZJX7FKy43iM2IgddUkDVJR5vJr/5OjFeCOfNog2ZLk/J8naLQNB9r5K0
gc4aWV+N2QXzYNNva/9QcvC7sijn1wYP4WVJMovanC0ShxHfsFyy9ZAO1yg2X01SrLF4vdfyRCuL
qM2rJdVesQwpb5w784rjG0hFRy70Yr4OQyZoPNgV9klFU9s4cUk3Iyk1KSO7OClswCsXjwqCMsVf
beUBof9Abz4gMRiPRGH9pYUwY1RjzygL4NvJHj0pHNdmg7aapcKhZZSiPYh8KzrPEvlSEaVU+SfT
zmqolW1FJF/d+tmHCDhHhdlMXmUZajGPaBOGwInN88XXKH/56plF4bpwxJoHSbcvzbFGCvj0xRdq
tWAkLbTJt6B7bj51UfNnT/IYTWJa6L28jRgrfwfr7hkWJ/hyIyv5WNx/rCgRJv6g8PsGxuqRI1HY
dC4LkNDjXHYSslOa6WJ20IlJaHJnrrvkAnbKhK4h0EHIen/6hmzAgzDkrhc+zWupDdfAmUydONZK
f+N9OCV0vUwTKmQwjDFxAPSpRY2rY+XKYomQFX9SZbWQM3HqDZFLkeK3VQtUECNfnwUyM9ld2gqr
GmYvmehHzkT4D9XXM+Cl8MBzx4tEepiZOMODttgWl5rRtc9ocfqAvbDCWI0xV048HF7i2uQvEZXN
0gr3oHk4sD8PZBFmBl4mpZMeTMT1tPBcSHqBIS6PYFePvaS2yOv+uYqRD0UE4G3hnSLG0oIMMAap
vELS+6AuYRAVeiIJAtjJW99vQ7cjdY1B3Nmi20lH61HpMGwVCiDi4Sp7QHXns0ii/sSbYUYhZHyW
d+aySucinzqOLVUPxnlukDbDHnuEKL5+hbyAUjDJLWTTc4N3fcPygunQR5nyqcw7xZerLFfL4TYJ
ekvIwMHHWNwor+P2UmaA95ebHCQutt0asy/oq5CBU1MZcnFa98CJo9bBOZOsWV/kyrksHyIR5IQ4
fyzY6wRd8FaXjzQwQL+khF7p4NeWxrVADFDN78Mo9eAq6jsZh+o4fjWKQ1UfIw7/d8cJsUG3+xZ5
gn1530nMpW6P8PIynw16Cy+Wi3TfV5CzzHuSpHTH7qoZ5UsC6GOFBx0kL8/uEWJVzzpI/CPJpUem
zZVFiWgWFq2VuPFOthi5bOgR5IcTEkPgBICRizNSnZX4dNPMwFtIbFOtn49DgF+ThChl3adHDTo6
sh1rnswVila1B9FENTBkr3h2buhm5keZ0uDKzbY+SOT5vUp0NZthWh4ArKKsoz9MESax8W6xl9So
64dbWPxqoOyWwpqtKiLqkyX9xl7aXiCLfOeyFZYezU3nqeW3u7UkzJjbQaOZwddOFK/+uKEd+ji8
jDRUksyZTC1KqT3i3SHg14G4MqI6eo6IBiSK5Y8zmSFwkKLSmFk0L/VY8v26MBMAlUm5dmZ37GBE
haZgisp3nBfvbSjCZzHGPKdxUwLuJRm8aenmxX1/5fWiyd/alrNSpFWm+N0ojMWSnplWhQGw+uon
iDTFwLIQoWFbOp7f9cxWhQrExPdoCvZoOQBieSik/SZauQkQPkRrWpzz8/aETj1GVE0ucTgB1Kxf
a9zdn8HPzXEG+JjEfIKhXTqG9+z7HSnQFpUWVP1oiwmVS85/tqMVCRDY9NnPf4aWrDg3lZSQ4BEU
4m7qfqXyCOoilXPC7jOgl5Y59XAvX9hLiFe7iae9tONNqbTQ0Ci7+TbDd8e1v6apMQzv6XM7hbw/
z+f9BckbxkM0OfrGmx+neqWsnifG+MC5xiUwL+QvXiO3esw7t/6CjgD7DrTJHTIZX07q92z6NIvL
1KvJRGc5RfB0M/LahIrgIRT3htJau9nBISMyvtf4EeEniNh6HX0kv2arygQxzsqtpLz3YNMjHgmR
m0a1aOVrljTvu5oJNtOhCtCe8gTtLRtFFJ+/yMpbJ3obpCAFJdWmdNtof0vBN9dZFtmlOVy9Y4q2
KX9m5MGqf8HtqhBUOFymQo51Hj/79rMCej/r9qSfMCKf0JZeRckgFdR9PgBwr/uqRalk3uJ7k4TD
9RwOAlGmrGZR6Cu3BskGH8bu8OYthSIMJ9me3EAnrlLTHJ4Qu4/kwGrtWfdb2ZWDV+J5UlHXjjWS
7rv73BJHpR5lrHQFjigdjUF9eTmJWaVZmi+2ehMnJkIsaJN+8OSZ/WCySlvy3J7pgCqhe+bnipng
NyVyOtzCH9EKnbZjZAM1sa6GaQYXxcKWq+VaCq5s0kSbv3m4sULcCw9RkRVpHQ1y17EOT6ER8ahW
MfkSD90cHSlQrSKdlQ3ycizPCUw6tL/sTF2B+RQNqiuL2Lvp+HC0JUs/4KGnuOz9YuHKPXaJz3Lx
AmdsyOFssnFIGMC+z96AngTnxui6ZQd6PW0+DtrA6YhwjmPmQCQ/IWMltsBRdu3SKqSjeh4Pkl8/
j1VyisGgbHOQcsVG4rw1aftgv+W56SjZmtaYTTRy+xbOJxFGXmiMke38vecJTB2yCfJNfxjNjC0F
hTd1ArgB3jcyGY/aPI7il5cqMFQhyq010m1Fpt0fCpxbj05gwKcAsYlgbWmiLay3oOUbuaCyx0oc
caYlGMSGlvm5YLEZoUKdUjZOXRmvLb5GvXGNHURJikEZzmObJ+MF2dOcsVioRfxUJSLdUrH/KCJe
3JHK0A9DQ03zGf50rhc9Hw6yLerciBySdhuPMm8e1BG08wOpMVQBy99fnz9becC0vv+nSWe5ZbZk
JaES8ux5i/V/QL8zwL5Kmat4+DB4BXaYL76VvOwIgZxFZtIFZ9czUO7nAIMAnHI71Nla3vnBQyfT
+RCo5OT+UN5IDiCp36/QHDDnrujKfYJpXWMg6DfRpvfHwBbue9I3fYVOYCm1arWMtc74gYf8qX8o
LTnQFagfCXD1iXibtGIiNlRF3duvS69sMm7I6qPTD8JiMPGi5LCm7x2cGfqXFGK01l+ow0o5OBBd
7qOnBk5F9d9sCnHh/PfwOB2IAf0cBlxpykQjSKmK3xWRiSa6LHL7eskSud0Surcc0tZ0n2CuifSv
QLUbwInjAxmvmtN2F6vckunoq20r8nBImDpeTmCvkPQqOOZXQuRsuksjCfJmbAun3ST8qI4dPq9B
G2ceo3vnSuKLBC9KscHhfT/ssKxnsiP7UBy04nx97cSK7rBFBLmAhLZ3A+dy9PF52JHTx2lwGJxX
09k2geyuXZegDllZyr0sGfUCbsHl8ZGSu/K2ZRuf85GbJncl6zyRlW0CNYeps65BVdkkQE6ccLGr
pFZ7pWR9VVWhD8DETYtlYJnjoZqAs51cRm8ym8s6YpYCUS14gkM0iyngGddxnNpVNfZ62exTt0+4
IwQMy2I6apZysWTmiJLuwVW37Wmj5M+f2lJCi6gc6YyjQHBXwGFwmxzJwYqvwGZDOdHysWggnfXC
QfB2P9MAp2M0iwEOCl5ox773vI7HLgaHbnIKTbtjZMmDszl07RiXbPV86c5pE3e9A8zzjnRF3b/y
HW7uGRS4MtZI485/d983lFQZZ0D0P2tnWNCpdytIg2mAWUU/yYZsOjNpaduRUAc4EtjFSi2AMEPX
0ZwwSOfKT3Sr7tIlp3X7Pnd7rbuGsIs7cjAnE6PpWPfgnsMJnZ2499S8OqM1+nYg+vGd/CbJ6ToB
9QsUBVQN4XOk6U601eMuR3u0/U7lXD/sweJNrlICNqQNktJ8EdQNlQsi3dYSFv2+AOLOLdeA4nQO
Eho50l6Ls6sMEwGwDiwTOQCTvATfg5klnzyJBBvKuftqplKztPaqQDKtVvAJ2N3h9kMhyebiLnSX
5DMrtJ2pAvhB8uHQLBi+EHQCFRdokXAc1xO1q7xkTTJm5Exsy9dNAhtdDn+ma8afUcbQK2dHX9/g
u4ryLdYNzc3rAhQp0lYwy5dJwJbOnVsmTpd9xQUP0iKxldh+4loQJhEGIKTmrI1rsbu1s49Dtn3O
bFMvm39nFPyEE9bhysQ0DK2xnCZV7dV3oXxqwfL8qhTgBapfJoJZh1yo1qNNTi+5vVrnObQDIAXO
W/ADG7yKs0QX0LeklZ/F/c/KEeyYjQJsnM0MJ9TSjkB3/yD3luLEiaYDX0l2ag5Ikv5SdfOJ2Co1
pQ5n74w0phiq17uJQzP2Ir8ptVn3MaRGRpMGJ1mu+1/NYSJ7skXIgctiQtUZOFfWpBighZxoOkDx
gSO7AQ25jHEnHpLg+5CmTPzldXVbHfMLTQFluXheM+ezfbVCPvaH2J7DKXWMAZFd0Xeb5DaiCFhp
9O6TQhcw4MXAhByfm8OlQEPmSUki4HmbS25Fk9tHAKHbztrIAhDF+MVXmwOIOwZKtxQbQ4gyTikX
U1kKVjeQ+40r8NXNJpU6M4JeeJgMFHuq1EfjSJdSmu7a6lmnfDmH9UH05nLMt6nP3Lk9DXMMmqD8
9RpbAIUeBf8CN+IjmidFBZlCY0fxw/0iUT/AvYMwy10Y/NNMr/O2J4FwhSBv5egSd3BESwpQOWLR
gYIRAwIM/6RPb6FynaTu7dfJw7cemjOOQK2v9UgRg4Ow6SFnFM9pdX2B1HTPzCF8LLbmAVFoD3f8
PGlkgRjAmg/b5Wllz1dUTKS4FQEOxXtBVu8rR6oKjYy8rqWJldl00rvuP1LevjwibY+uhOawiSAB
jtjyQP3Sx3ljpYVqz59RoESLBMhlMqNMbUJGp05nxe7G9myD+9v2ewZP7+TGYIE68MRpiM6DUf4A
z+mRYrPg7jH04Siyu+HvjuJqNZdbGvb1/fNEuWbytrP2pADyV8pMz75PSTBgKTB/VKkZfhJYLAC3
MsiJL49TG9FyVeBX522pueNXU0+NfPQD85WBBPQWaJldUW1OV4ndpE1U88p4sExRXk6zrBFuu9tt
MgWpFhJjMb3VzaHukye8djCIsmw3RvsdCh9/csxyJDW0zcAEqY7Nn+7njezpqRtZ2rKJS6J/Leg6
fkujMRGVB3cegsRPgsi6dSUChjyO/A38mub7oHAMemBA9qxGSJSbQWZ/7r1H5k+KOxv9boCVhWd/
vM5y4NHonuLP8BGtKZmTtXRek/h+PSH93CH6+cMAIHgI3XvAV7WjnORQnE36HF7XTjjyDXIki3ef
MDn8+6o8y84z5mlpPGQ3QrXh9yILl+cyrREDS5RFZV5Lnga6vJJ7+2TDGOTdZ36wnL3B508u/oGK
j0QBUot1er1IrNEVu9t1Svq+c6NJzxJZleZFdHTo+cETrF6BsLEpyHVdw8Z4yx2GLRLNft1nZXbJ
ala+yfI8lLJ6tITJc2sVelASiO1++rBfZg4HimT0ZVF4yHYRgvkBAq4LexipUjHb9D2DNp6ND4+v
D8V8k7VXjwnw202phEmkqBEwOtKxhhSIgnhdksQQLv5NSfZ2IrzvN8yBfRP2RH/Co7ugTsuRE2q2
l0+w2USyoO7YAhI2SxxzAthl72gQxa+3gbsNsIdkA+wByz5Ij2yDuUPbi7tnwYc24/Mib2mkvlFA
nUp9fHzLZtIYP8Y+fARB+vr/+9g1GCXbPadPi+ZPTSjQHux894stfa6qTX+/kE+MxA0x3aLBM/Tn
7IVV0Rw/6tA4bAN9hxStcsu4DqB7e3mLmsu3jG0AxzTnIKVSUTk5stz/h4CGYxTbsZly5pixVYt+
OpSZ59qANmhzhChEIIsJgiK3vggBh/KLu08BDJgOkpXcmklTNU7bvYqfiJlUONzVEvFnQtFHgS9k
m2G1zNwAGuErkzWDbo9uE1opqBCevx6xz2V2jfAtDpqE+gbfnqA8UXs468eCh436Ogs6RiOnuvAS
UJpPhl4HXNxkB2oEMzvgBXYBPlu/3iiMHQhUuqMEmcgearlHWAs07ylgkWeBnVMNtADVJut2Ogp+
2pudGj+fLpRL94LXJKPXi68azkPjEk6qMzE2tQIViaBFLKKjojLByg4nzQdnU8oC78fiyBmPgvLd
gs/fz+VdIyS2b3pZBDGdTv/AjZnufLuhw4SLSQTA1NEasp0WV7pmYe1d6Nr7otgnP1Lu7un/vDWL
1mnCyLNsNrdP1LqcN+M5G/6ZSlZUmpLKC2Pw56cgLpGD1IbZgQXHpry5HOyqARMBUDMf/e7g/W6B
M95A8+kpyuu8YavodpaDS8oJWXvaEg4nGYxjUqe1aMe4mZmg7S1rK8jThT2ZK2hq2hs0ZJ3d7eda
6HYmxbh3BYxXLdeYtPFl7mG00pGnLDqusQzU17AFCAS523T5HBxcZ3ZyM1QsJG/kd0XAoNYEsQee
PPyB9TnLtdByv2WVCLA+17MG5ZlEXS0oSsUjD09eCiKViu2QajBB/oKW5/mrsgJaUrNTHlrz4jMr
7G5Uq1blapGg01NLiBaSabXW1TlEP/2rmVPtAgXrs/ZdCHxsHz/6lslb4PuGpBLEsGUo1n3Awozy
Al7KEzPsy+yOqNaUJ14Eb5Svw/CjpdPPzOXftZMg3i2STXK+e7PhBNcPFR05NtklLm2qehfrhr2v
ddRIWdk9mKUmYlTrhlX8QCR0NjhT+qwBaDM8XlEMvNA8w3rjeMKZvOrzGPhyfMexD/nouctfOh7X
7L0a8uiOZsr9aPNT3zjV041xHSYg5gvJZIYu4rInU1+gB3/xtGfp9idb2UNbJ0TOr2SzaenSSliB
j4rXxIA3CSzMTsmlms44sKNIUwdILqBkNXqSYW78dhiSM81hdzls+au/UZDqHvTlHJT0luRsdwbZ
ilPrNxSBHXUEz6gQ6UK6mhU7Bv7LQeSyIIo66g6uZPn9ngp6zLe2BX9g+FoH2KCb0MJsBaQG3UXF
ukb6wPUJjHPLVqjkAVu0jZ3elkZwXCttEQeAIUjBhM9BJ+/vS2V5Tu1/jd2oNVT5Z8iEzBBLEQAC
Y2l9eJVyohQBSQeLd7X7JOwdweoPjo27nf173MTTahTveyIHqYXmrFQIt/EUcGoUNr8pNFJcMzIC
DnWavnidrreqhOv9BOQ1OWXAalYUjit+YfNYIxKM7CnelL9MMyImA/EZ2sB0xO50mR87u5NZfVdC
U9X4Q6rNFIINx/fhM4sFirOYQJQmD6dD9YPmFP9yQJeyy9X0Lm/ULhtLMiyjSBkW/Dk6I8zSzktb
wv5ekAS82lfuz4HaOgZHCAw8A6fC5wUWeRYOgUytSwfu5BlxdP3sMGhl4TWtoUEFtUFjxE0DyNix
3fNElyZEd382+i/ziZZxza7fr6DKjEZQ9llqrTKq1lv7fKkGRjIGMEa8KPdOAw2CfLGsUkg9UVMK
KI0r4Gzyjm451LLYZJ+mAv8xHCV0/wiDO5hLxsS70jIBqzxld9hABtp9Zx1RjPoUpYO6oO9dyXGT
y0fB90saXGsZBDT3BtMdU1tnG3dN8GGg8hO7ahCycC5GiHfP7vpvEzs7h3bplRWVFNTmmTbFl7I7
3bqadbNdjAmtC1SwjGGuOGT+4pj7RzfR4ZkVYEpyKXaK6jwyG+KlV2GlqTTkF08v6AvG4g8wWWAK
cgnX0ekJNBhQwUqrFYg9GYMkv5BlTyBQPMM4zLrx/PzrBZSz4tz1xmm9/yCzxCrt7kfg5t6Hf9Wx
dwbWtJQ9IJBaCYyMPZkGFTqVQTe1ByLKMq9CPyloTpOwA8v9JSbukzfKkSMhd4P0wchtWnPKSbXZ
MDgMZULaHvpm2bjoYZEWrAPTy3JfvpCc9yCweqBtcuid5J/WItNHsAeR4XMTrJEf5ve6VZ2Ff+s8
I65snVnP//egex0Ur6S7aSQpkf+ikFQqE3EFL8XjwkU6x8Detl/juQmc2f75uvi4zgDjY7SBEceT
3fHDPMZ3/vF/E9MOcO0hp/qLH2MTpAa38p7mdRYqTws0IrRcQgvbwRUuf/WYBgtHKnq4h21ySOit
br3AOJIVDzpuOKAMemw2LNqEBM+sKYxuJ2gqblpcwP++7VV6ryMxgtQ3xgehJKx6v6dnsA0d37Dl
g6Py0NYV4dLI1T4vnumgcyhxZlZzFeL3sjOjkry8cBnXWqn+mE/pfBOw04Jl4nxX3gSJKZOeaAfF
7Q8sV6zkqVNImzOivRFGwhPMeTvyO8RvuGhfEq5opMs7CxsvYdgEjMGIa+wzqydmECKOdX+Pbcsi
phZF0/9bJ3xuE7eK9HAJcNzgJdq0c0Kr6F4JnluMkE2OK8ZiYRMp6xMOjYCAWxYFIQQo4fC/3CMD
URtZtAoGYz8MsiUg/kDdPVzAMPTj+ecFR6shmMXHn3kpr5BRGekb3/rQeQZmI5fvJut8O2BoWduX
FdWDEQgf80wDk/aPpAr+kkfRBjFKzbkIiE/ArxRyNogEzXRTS34dKORgXsTof3lGWFmkgowwO4JO
f7CRTxqtkSVYwS7fQtZtwTUMyuN3iu9zP4VrIvfjfNp7O8PI1DYswtpkWE8C26ulIwU74zYLuB9t
sgiovfbgFkehdDESGmbbN2deexoR8ctnwiGf00FXk68byc9sGtCaMifB3faW6g1DCTzh0cSq6ZSZ
wYG5wMtoNpf3rV3xHJLwBEJmNW4MsvgPQIA4YdXnSee+DvjJ+/WbbK/4Lhj6xiQqgc3mIUxcwbCP
sG64HZz6ZLwpiLFjLdJI926p0dnDVJcvvQxz92B95G5HLOMxFLLJxlr8R8aviHO1WjIedCpNPVBV
VVXDVXSL/VDKlWzK2O6GLcB0yHQM2oJLHhIBlGNKS9imt/dVKOxOmB7bLkg21ebV41B3lssJMeqF
SykqSFARr29+dZfRNNKx7RatQtrbnhgEVqbUJtyFMFoBmAIWpSEH9xSteF8EJ0c1xYzs0x/YGsLg
vsbUwGxnthyLHVCVaRWOgpXFc50b5oMXy5ddMJA/19YjOIeEQvWyqvp4IqpkmOvC4Sqlz6yL29uR
oRn6BO35f8cyuwYKsY0vpyYy0SbfW30wufM8z5rxw0XyrONn0XCjx5ujYVXb23MOdqwheP2Y7Vxi
ayo//rcdjjYbBCDUtVEgTLyhCfi8AcFRYpd7LD9Lx13BroAX8iSBoG9wV8vw+APChwHnKMaf9UiQ
ubZ/HExUdvY+taseJpQjo7ONyyq57G9SrSOSe6eOWjTCzCd+SKgMMrqnjsDB03eHcYNtFYshLKhZ
t6OxA8rLBJfGjq7MkC6IqUqXbATqhoI9TW3JV/uf19aNHo1BpUAEeIItwv01nW7aoq51lJQ687Jn
Y9plIoUtAENj77lNWOcwwScLBgaEU8Ncrn+MwUixRgcWKdLW3RoQX8KiciY5pXdd6C4CRx8y1Exo
fv8xcjEZdhmSemu5tDkVKKDIETDNYAf3/jO4LOsi8iIHJlMVL3hrW8iN+l/5jBfu9JQjLiP/XSh5
1x+WsR2IydK9TJe+P2USMt424N3CYH65z8UEDvG8jU3O0U8eZzWHx76cwK3OQaZy6y2uaxdRt6pY
MO+geSBZue4KNkOG0LyxGGL4jEhmgwtAjiINw5Re84v4Mi+C/cm2JiZ1Wh9a4gWBSiCmo7qCZKHE
MN0STsaPR774wxAetT+igMHF61f0wIC0fAqpBBLVfX2ob81v8o2cG+6BM7KYJoN4shAFvQUMtqd1
klE8YZcyDemmp84QxisdpHt7S32In4c92eZnC273sjSyouElBlegkMh9s9Hpgc9sUxvS+G77kvJT
96NCq9AzcCH3HPh3EuNVvTxhEXpIM7ghB59tflI8UaEXbGgimhxo5BcnHNy77OnlTpovWJDjbZTv
K76oVEO5ksj+NUpVq8V8OuvwRFftI1kkpPCoVOfZr95L0S1nWXS9pwqZGwuqzSgznaGjgHczLgkt
gqmznUhxSlyVQ8voRndsCgkmXPFdbptA4iO/DI+up2LDo/q4+2xPgrPdCmphVT+TeUV1JyMRX4Ht
/4XhoBqwT1pas801F3peSWbPez/jJIt+a1WBlUgm8WCyz0O0auQKhQesC2vsYBTH9pOK0Mu7LFy8
dyMHqQcV+XOIFREeuAysHeJ9Qvy59gAbH0MGGNHAC+5/l/fDnGpW8s1A7Y91/hRoqsrJ+rrhkOhX
AmFZ9qtlHaBayPtbmGPBo1SWyCiEraIAp4O708LVwXiK9jsEE7paQxDL/r5exKX8MUTBtcG0Knyy
SlULBkYfp6mc38zhQBsF32XoW89uoZg9wG6t6BpWJ0El7qgBkmKupjD9XmcqzrSdIh9aInb33+T2
C3eYnxb5KJQ2c/S3eGOkprUq6G4GQ+hLggA+EhAOn9wBsWRD+YJJJ/ZF5f4zxQO4t7Ry+SA2sxYD
X8q+zxPodLjQYBN3dqppq79dYKruazHxAasDoKlfjCbXrOOrKH8Ju5r1AF3JAGTaCc6+P3Jgbp5Z
bEFipMdAR9nF1Qibo8+wYqhvFXb1L1Ozza+7sxj14Vy5e2mY1HgYf9aGu6L2zWUPnqFQ07kR23qG
NbZvpXHgpUcdi0N4HBH5KBzXgWRIWC3IydUAl33/q6d7EbITMZNGWfJ+d0NIPkkMelNE2/NaAZDo
VSreHXX9rtmm1rs/QUr65TaX2EDU7WunQEaG9IZWIfNvp7eUmRWgCBfpwdfijjP7MmPrCoDWZpnl
OYiX0xJcsfMREHGz2H1GNEJrf8uyrNsCx9UhNnNCbmGO7rB7yATJEVVeavG49LQ70084wTqrXyCd
h0HBsN/+PfJVfj4ODiCQYz/fe1T1w4W3UnAxBrOmnL7x2rN5QFh2YOXlDSSgeMcshE/OhJbXHLQs
89ESOMUJjROMYMCdhkGE5O8phILoOgyRvyLFz3Axu9kSXBLT+l/ECV/Q4Wa700itcc6ULllSxnU6
4JOz2Zb/b/EFFbWxTm6c/buG9yi1lpjgXQpTyKgsRf2Igv8lL3lcpzCBQSp6DYcSRqqIvrlhqYng
D4FWuBmMl73XUYaQDWz3RhxDD42FXD+gfKReiMDm4MuA4C0Riw8qOIQID8Ctw8yfS/zzFBMVM0Vd
EQb6bnaWTpsixaI5n652JplkRddFnJLuikcwRBMvp2TFGzsOFZChYGcqBG4E1Ue3lTFo534mvuHk
QpGdiZEUs279/dn1+RQMTBDJGyFluNm5eTsGJEuzAJX+KL+fS3XanoDFQOd+iE2rFQzBX7YOyTVG
7/zhTn932Y/SC6yd/9gjYBTU9xLA9My+kgjW2O+J473AVfsIdZ2C85UuxcJC72uB9OyFf2XtDZq3
jGqc/u9/mu+4RY599bEqCyqaDQY7N3KjOSRWW7szDyjUB0kUNzEhccShR+jQWphtjfJcwVlpKw7r
dw7hNASUUWz8Tyc8jQPiitYGvQtP+T4avs/dGZcuh66haQixREJOT3A3tkEc4AGeoNZWO5dvcQFW
QkARtgLlZ/aRzL17Y+cg7fiYLcP5BK567I/c5mnDNc0Hh13gRp9CHUYauVtQUv6hygyedjcZbJk4
CRz6bv6JU6oST9TyGLjVihkJOADJCA1YBzNNqUGGpqPqmffIO4ZrzVxmKiOw4i2z0VN6H5EzGbLZ
z+gAHxL24pbobpqQDyjnqIuoSqQjnFrX+CyfwFbg3040o1WSLH3Pwn6uXEhr2CeSo0Gg6qgE9lYM
ujfAbTe1CyZ/8N3tK1LQO4WmHpghGNl+/l3QuDz/dk5tjFpgfinczVhd7Rk3m2Of6qwFXu8KTiTQ
8wtF/2q2APCuFzSnSmCMyedgXcg9BXAMBxepqPg/zEacWX8OFf+Wzt0ahvk0+4CNK/euwJuC/Jc+
p73mjmRCdS7QRsuDFjIqBIeHRWeC59C/7B1Z2bP1gsTc9eU0koXX16hqT/fuhZCnVAF1I3p1UGwr
dJD4UMIYQOMhk2QxmdF92Id6ORaOCcFDRYWC83xNH5oDkkSRgFu+RPPRHGOf1KLi1Qx88Y4UnmCz
3+axSTO3VCfg528hWetDBQYbf5uTzEAsCLGCatlCCtLkTRtEsKG1ELlh3yehFEaZUBHeatmr3SD+
D1okpX1l85Ag52vWfAo+KqRLytCLiynh2vOyP1RvnGQpUZP5vWL0bbLs29v0nBEl0+/FSegjZ1/z
A1GAOqbsFvmBtK2xlk4Ct+Fj1KJFUwUU5UVSsdRk978C7p7dhik/FhObmbMEPdvrdCj2zSJdfeBH
RtxnupGxxj6Qym5XE/DCkRn+BIBZIBlW7bCn2e2g/h01V+G35M1SymAUFHYzBRqYOuqD+6s4shyQ
0dhqzSlDd4lgQCNyqQtuDwhouVbugyt4m6r83ouJkHAS7P7+pH11hUQNxme9BpPeZkaWfZ+Xk8mb
iYa+XVKjpRBv6In9KF5zCTOMQQxld4jSJ7remxwFwV+Ipv3WBjjIEambRqqJlil6NAs8cscrd0YD
GYqBYuxwqxSbb3vRMw1KVHNytBQ9j+fCkUYmQzeIpVhLTFBxHbXOQxfoh2A8pbJ1QLexieXwJ8BI
y1JNeyH+DP2AW8v4xwpNemLduI3rns1p2YPCdl5s2RRwCk02tXIJU4yGHe5HVk0OhqGOYA+0c3+9
/qC5T5uIBo/7a3wusUlajW6IxeZLg4cIPqq0RwsG2dQDrp4JJbGtvdLNiNYqBBD5PTWIjuxzi04Y
Y8tQAlNgDxNOOd6pdfqW7ljkfwLYbzEgv4x/78TrgBS9c813+91X0P7vLMWmp8O217KN5eo9ID8o
fwEsJNa2meLYJd/siyroAeZQlYeZiCPbz53UZvRZadesNSKwFr9oy8WAr8yUvucTEgVwLJlt4jCl
XbtAMUeqbLl5HMKS1IZI9mvkMg+uT4X6ttiL/TBxO6SuGj57eNUqd05TnAMFNGscLSk8MOQVTrXw
vcpBDpK5Wtjm0SxOqzBjnP6A8pBb0rfAnN4S/8JRMuOJ6Ls6tNTStIrV2oMBvT/Pxc+wua6IfMgV
HNAzlV1ZH+8Y42zeFMjCTsGRPKIZ3SMGQASPI8EmUVYqMnszTxGTmc63Ep7r294PtNOlAlCxRD0g
TEG2N7dDW6apQp8+C5ipm0HCHuzjWfgv69mn3k4TlkM2dY9mscM9nADf2LCLWAbvRCaR0uGqdacT
Nay8p1Xr1/xyN2nIZKqgZa9E/VZ33J0oNq+Y9lHaKxF/FQs977z5tBkEfmCaIEbhDNPlSJGuBWB0
2bJtPtdFM+78UkaJg8NvTwwMYhqOdyU9muVLO8ABFkLTdvWEr2gEBdxRb0cCaNT5nwtbLILErcVe
A4aWijQ+m1Ks+SBtn3ffiNs9gldPm4S7BrlfwW6kE7I/7o204lb7ozEfPKLvRcrGOuX6U3Kx7Nhc
FTtN2G8w+EmWEgebq+XFeNW/SusZAh7ez26KL3aYOml6EsKWfceyQA/NjsXMytNGo28F2I6ywfc2
F2izT/m6l5nQ9fOKcGp2KWY0lze2qDyolOfvQZUQ0jfn9croVa3FUm1g6gYSFwqQRaJ3bp3REnDw
FiUkBHPxakBKlGdXFPvvOJIjT0ColVgM3zpQKqn8icLOmBtzix7dKw8rnp1ZT8YtgO+59z68i6Rt
pA29lRi2yDtLNfReDxI7VNPIv1OiEd4VmbTqxOYdF8AkPbGvVaAilTBbi1MW07zZUms6a9Dk38FF
IL0RKhgipY05RTETLr0HTXw1QN2lTaCswi7WJ9nWH+dhzS5rxLvuitWIhfSnTmv23UEibU14crkh
SoNuUcNesx6GAsGcuFpenUva0qNJ7ZAX2qLhuDwSunTxm4lhQ2WHk4AOCxM6+xAu1HnePFUOR27F
PSjet9zG/NZ3VZ/dVo73RL5EZb9KFaKODOheJu0sl5Zzl5FGtQtrbpchbcQEKZH2Z4jnZasT23tF
uJ99skT6Hqg5nFYgkRHr8B6CgWGceY/Djux8eOboprvwLIiQ2JAa9jQS6mYpUWzu4wBIPYiw77Ub
2U7Vt+g8ul2X64CzKlwKo0CVqWManZz8gwTz6JUXiPIaMB0fflhA75q2HfhzNBeUbVZyMmXOdpGW
4HruAkdoWpG2DPxXHmTQRWRJEK0F1tQdyo5n0W0qkGfOcpNnOULWscO/bog0XYBrX5S2WjusvmIc
PWeIqK3YK/FtRzg5c03fhVXiNMcCKoiKPJsLpRq8n1OBSMCPJZzIIKF15PC71SUAxBDEMfmFllNi
yNYXBvr7LyME0A3JDZOwrbuaUhlxTLcut8rE0DFi/+NaMCR/LHByYSQTupGOnq5hgDv0Gi/Dzqwn
HduPexYa7bfR8mIM1P1R2XCsQ0qDBPoHYFPl6/iy+0FpwoQcUByitP9pCiQFR0+gEBhnWPUNFTdz
LVUI9eKxmtkCNgSnd59o+59eVXuMPfq5+YBQM1fGfWbbVKrTzrv02KLzfHy5IoSxDFR0UiylIKmn
KZ4zMIoj2rHhT2iEJFMKLlatxtl5S30hDragpkjvFNDezmPJzjTx+IHVgaij1LXvIms9qrlvknPW
8pqvYKmgmE+cT2kthMXKN0MAQeyFF9VYIKReQwykTN8qE6XeNVJmRRDxRvne04Uf5sCt/GZefbIP
zPdMYVFlmJBScmsk4w7FsacERtbZgreKEH7iAUtF57U1Z7Cz1Z908e+owySXqmkR6dJfu6dXYz3R
iR1U4xArC5cnKMb1CHPokhxdXldzktyBJyZ6zXma7yclK3mXe0y7GLqNYX0uFmA0XPGLyolmoqcV
OTueddSGrJ4zqRStVbPcpVH17MLGy3kNSHAVzHJ0zvhJDp39cCKp+JVaLl9SM/p3eRvpZtaCXaQd
hxAB6S8Rb7exsePt9SaCoJ3e0s3dtX1aUybY/3FeaufD08Rvm9H2772XudTsijQsPaPrl7XzdyWI
4WuqYkSFj+WsHTavn1Il63ZRDQ/afpjdyH+H6F5PC1p7PhgBBFL3z95zlncr0P759ktcZ4zescP7
WcqrKI7hFWgE4bPKIFlT6uRu23BqJyvjhdxOpPdBECxnKVxgmpc5nYK6/RF9gAftvp76cZ6kSkty
PiRkMkmznyxjB0DWSGLAvdtsLH44d7CiXRBu62j4OM9kRncbe9qvTjeiJ+fFmTGoA1/KlX0pNujR
tHbdf7aio44Qqla2i+4Z8Hv43TzITfCtnIrzYsuHEr0Nc/LROsO9IqOASpZu4yE8t60TaHVrazQm
gJ+5RdXeAz0QYEli9xINKz6d546UiBBsCQQw+G1yOpAwLmjUVEf0l70Wm1chbqr+rUBAdwGw7hk+
z92sNNbOT4HMkuqB+Am6udl3EcrUSHMhtlFJW5myYP1zOVCDAItzTpRAfVZ7xYQvmP9tmN0E5Y2U
3jAHkVSG7msCzp26N9Jm3f52FtjvoRU4XQ14PcfQ4kcaivfdkhucTC+diXek8Slutmtjxf1cMrLg
wHc5gSvTZbKTgqgmQu1DpJ+6Zi6cQpG3+DF7p9QLQDnuBk5M1Rx7hMvDqGAGEYB75+x5zfRhTI8b
zPi32esv46ZJOf4D7sQcu3saAnCZo23SmWZBw9rlr2Pu/AfonQT/bAczwRGJyjQFmREY0JYBSGaA
QI38RUZk0gZP/T/gdgQa0pYFJIDpsxDbyyJDiWO8DCmKaKOeeYHkS/SBk629GYOmRHM0Zmg/g/ap
XsJMqKudgXozlq/QVDt92fakvuDhqzx+e53x8D66o/p1MC5A/l9DR6C/6PDXn87R8XosMwMdW3iP
cfkF4fnI6IsJHYTsiTxaPRpxrTyv53a4GliRT3xRdKxM6wEl6JPCNBZdWcWJ+kZ7zYhbF1pNOHH0
zrocItvbN+1/wo/r7jEsOu/n76rEu9EYZAWc3CiWVh62cad5+G5sSA8a+6/RGkQNWKHvxmwSLiMU
s5tDCWvfeS3SmYFj0rd026jmEyPk5biSP6sJiFPEZK/el3myFTiiFY0sP3nkPMOplBWRD8Ivrez8
QcI4GpVmTCuGrsx6ALSagwYmpXOP4dS9e0GM3giUNmmW74hO2mWwH72axXU4UZf0Uv0KnDMOczLx
2t1bGw+F39HCjzzqmvafcmtjyRKa8MNhpqW+m5S+PA6FMYc4drPY0qnx1bYtimwTvFd+5BDk9Oy2
2keoYDTSS0kmltg/G9OS1NGPdVH3tcwP+jYDMqFVsEn4Ww5u9Lv7pU900TomcPnChnH5U7TJHt0X
1K/M8gPf5LP4H6VE95rBgj6RDapMwztvOQ6C6MXGebPyUntCQXQfn1e2TTI41UeoSaUfaZqDUe9x
RFDTNjqGx4HMni+HDFFATH2NeoVT09nyBOvyUNwjOt0FxieRS/1mjDMPgP38WCh6Yl3A/NXj9Tfx
/XcSmI/3t7UIt+MUy0woYnNHtKgRy8B60/ZfrHdRJRJmLM24QGO0LFfVH9WY8eOzkenTUXGVXUh0
sXMN56/uiCC07+C/ggkAF0lgcKlh7v+SlkKtdi1YfFYRUdE0LiifJAqIB6uqgTG22iNtgEdSWYzB
P4kjgi3xVxTNk1EiTzrMjyvl9MziP6SQ6C4UoBWAFcKgRzp1GtKeVPU4QYiKeL/yumL+Mac6EtOy
dVbov2Ui03EVD4rC1VeE5gd730jpjsnKnvrfQk0gtqZJoKYU44YxP5jmmKRX/AWMv52MUXOzHk+U
WjA6e6oDxKMRxU/akqvl7Rg6JLcQM8yxNMRXdkqgY93Oarc24+O8oaq5bJm7cQAyC9SC5iX2a8d1
t3BFApOtSD1Cyd7IM+e1S3kMvgSimoJ1JdSQKxVPnpGJGpUhT1CsfZ4PxL5FagWGd2mVMa5dvlAL
mgxrYZKaDzN1/hCpW35yxZ5vcANYbjk0cpJOyQrP3eTGQtDFBM6emWLtu/YIiW28xVwAQCFebh9G
Fev4TIdGSPKlJmpnAqe197z1hiIFcCpjq3FoLg2RaoIDyHrUHtnlwhYGm4SHBqDdmUHbxMvfi0al
D0WZ9reRWk5xpY7d2SE6nUdbDDnEQHeF0V1GiJrfmJMm95PrCNErWeAW8usqHFKbvhv1B0C0OoWS
4ZvRgta8ja1RYqBf1m4EpcMMbmi5CXhMc152EhIVgi/urlKrGupyd6Gf8kN7v6xj/s+q1mBrNZAe
2/Gss85KNy/eL4NuvRG4cJP1s+L51whQr6vYurPmj+ri1U9eTZ1UCp1yk8LWGdLHKJVguNxRv73J
9YcsNju0EqnMxALKw7HxgEf5Dml2TWdwxcCtY8S6OZDSO4fHY8FufySltdNm7BQTlWPrXfEjgA6l
KqeW655LB7EfpRz4Xgmi8EucmO8FIThJLEy9q1vdF9v+khWCkxoIzU3eNf9E14MIDYQKltV8gO/1
itaNj5saCdPQbrHDT4y26dFDgcMUVz++kLtGkfI23vndWhMYpYEg8MR162g5QnKHeAgnRkuStCsn
7sSQ70AfT1yzIKEKx+17GQyLg6X55JIXtsA9KFMT7EQXymAwaBTBAJeIOpnabbfHkGJPl6b/dCXM
4OSHyhO14jfvIk54vOfeuDncPb1Uh3B1QNgZPUu5uyots2tlIseqTpQEgZrX/BaPaPUe4JjbS42d
Ntci911/7bkmnEHw2QRd1eMjNlBbkQFcHcnbp15HAKk884bP9F1KbTqLyVbPwBuNq0dwjA/ybPS3
B127d8+JhtBq4qX95/0nHEnfUlwx1nOWSqMMmeQYj1XS2XtXbyaHEKX5R/Y6KPoBZuaFihkltCIp
zNGRHR3+YfPPqfH2qk30gGONw3BnmM3lRmYQoD7yyr2u5sNKz1Ok+MyJOGy7hYpfE4cOKsbaU383
lk3ru86ExYlSAoHkQPdibd4x7kdrq7xiSbHJ6BBGhZdHcoRHyhfygCGd8BnMPFW7d54mK6oVA6Yk
RraqGnxqEQ0VbxA5EHvyqOvOJxnyA+lgqpEdypFz9FVPmALvHK6ATijsA2twoPp4CEJ0b8XLojlf
TMVqY7JA4L8AgxzF7IcngA8ELCmY5B3LC9+biu4c7p9c5Ih7d+R1HTj6G/Dt+rWNRHosgrO/4ZCh
jIIzYT0K1HTozTFtNFphxmMbenfcyLQH/uussM9vsYzTwc4GU67s2a75kfwX8lpB/1aldp8p9qpj
MA6PXXltvu+dLkomuz1Yb3r2MF6OqFdfoZ2ou3iybYmSQIf9k/W4Hf9Xkk4HWHkvaKU/JpZm5P8U
uIqwBETzhx5boLxJqM1ylJ1bb15tKjKI9jm69KbrXgO2fXc+BvPeWeaL4FPf6D8yEqfwXqokR/o5
jOsOCEJcrAehVB4XH/oztd8g6a/VNhYwI1xKq1koVuU60f2sPM6st2Y23xe9MbQmb/qO/xSD5F0M
LN2N+H1kb2MQOvH05rmXhLAQy78YfN7fzhFh2pc0j/XNrqVCYmHjTfZJ90BK3LYThVog5sPn8q4P
QNeGG/6AV+tkZcpzW+zgMFhb2UuGSELCxufJ+fGeibfhD+WKc/h02wtJCSULgKWuXyhv5KNjuEon
UVL+B6iycOzonMn0U5WkfyqP1z0aXrxyJ1UyvNNaR+dUQZkX/q+psCXlJ+gSyiCPorhoGKWzV37v
9MngxMxeXyC6nsBCvCTa+fo4gEw+0XkTpTc0ifra4IP4J8sSScW8WIqtL6gEU3T924q2gTyLYDF6
FB01a0JQzRas84VzIdv2GZKFB86P3VMWueYGXUt0fhMBFVAa1rN/r87l0DFL9uDltDMd30au7P+p
EnBTLXT7U7rv5rP5cvIfBuLkEC5AlvcGEzk/ouIhMKnzPBUdR7ema2npILcc30NH8WkbM7txn0qG
0etE0i62JG768/JKPncVfRIp+2IB4o/yx6sU5TENgzswxlJlchs8kIoWg0MBb9JZ2uhcz3fugMn1
auMWIs1BNBb9A22WB56417nXJBgcVC52PidBfMZj28gJf6EOVzR9RRabMKbLjULSrN6MEzSzCUKK
HDwypx44eYq9qAYM9RxCdf7IYUY5ScBurhIi1E625ssBeMGLQ+o7aIXKP/Ul6SW47BPzZWGBzZN3
/EyaPclBfvvYtZjmbGIK75sSE1Rlm7hDkVC3A+ii+EJnLFfNIZpXxA7q0PQ1a3HXwyu5XmfKFQ91
EkLiy1k6W59ovbEeK9WNKOwK56/vP9ZqtVDGbRFY0kbt9KZJdLvai8LOy5l0Kg5ku4WUuxbHOMXL
qGf7CsRKJ4crku0KZq+d9pabOvgrePIIrgxg1HOch8LTg+WJpUA4hjhu/+d4Ay97vKSAXU7Yg0cJ
CuBbeg34GmzKPsxq23NNwNbk973PlWMCKxjd5Yydq2qQsgqo+VQ6apWoOFIfuSg5lBl2Esz/zx41
nlW2CMktz5yjhglTtOfUqdlqTOLTNtMyCOu3/+ua+vxaLo3g8371xa/QZit2Z1bdC4qMIxrD7ffu
xGX+mJdze+YT1A2i8QER7R6POQG13KjfdZWaL06R7xV2txiSxhL79UA6d+PHO33D3GWUdKY457n9
Jx06a6uk1D3Vi5Ar+YwN8fQDI6zIUoSPKxh0abDiyjeqzkF31HP9DQBdEPWCqqAPxP1iOH9ekaHK
Y1mZh33QxttXgG6J4j1b7fCVrtjDhXbxudSSr4dh5WLq1sGvSGN+pbfAy212rvvVPOdbal7Wbtgd
Zxrf/bY6X9eGvsS9F3Fuv2OwPs2fMbzcKH289o++b0+ZYc2FViuW2QrRS+AoNUJigzXLkg1YGTjm
GYQ3pMZBuMCNTEazIAcqw954bmGHWpOmPt2LdRn1+t/vQ1WAicmD4MSGZQ0nBsm0qmMF16s++0Zk
VI3Taea2J7N4F37v2BEM7pPdJn1HM5frYqAkYt44EFXT8Yt/36myemlaeWGko1IsROkAqJtBs+dH
/tmU0JxMM72S19lRiIctpfISYFJtm/jx/5ZV38NutjfJSl84+i01O1WQ7cbliH+zx5xWI3DgUWSM
X2JhWBAp1WaFhXwBpOTUl0U4H7+AbVOTY1H481Xtu1isaGm1nOJdxX8i6JTAplmejv90Q6rqRp3t
72wNhOtRFIE3XvPJ/7Qr4Dyi8WkOBikpYmbBb3F7KLOXhQ9pO42gsHcItM/FpySsAXXMVNAceiIu
tXEnejLNsfFsC/KxnBGlbYtE42MRa61q5yDs0FOdpJFklLdVGJhZ3EGdS86YvnzTpLk1Xh+rb0wj
ubD2FDiPSpwdYVhPts6j5u2nOP3FAKPkvbL97CPJM6N9HVaRv5F3u0bHtAVAKMgzb2iAei61yqvK
eVLkvz9kC8oRKT9rFDzqr3C0DsQ67FimWsZkrUvtZHHlAsmQzBeZ3thERts2yS62/tBiq1XaZ/M9
mepzVTREo9TblpyaneNyswl1/mwMqnE7lduHDRc4cvg9NKYaqIqpp1BPVYou/AB6kZF6SHG/vyC4
uEq4E9bsj2PAvmQ0D4XxLT3nEE2uoGnuk8wtL/kst22UFFo9y9R4Y6PbqjHo8CNcTw+ap5CIksx/
6pBQqa8Oola24l2zIUIsvc6CVI8tDCilY78nYnpsjI9yNAoOe3PXcvo59ex7VnGwxcWsrWejupl/
riTFEa2cVIXOmqvxo3smvnGsTZBHL6Jr58II+FG8HvNeOQrjaf+feKnKEf9CHjiKPFZ20qd9D2wE
rSi7WYBGvwc1Efp85h2ZAxnYQzQH9hI7RQ1GM7z+ye/fuN5/+lgtTogeVmuDG4v3RNEG7cvDs98e
XucrogterSG26Lw4dpybl8fLSeu3FeNtKHCMhp0IE9pWjtmut1iR47Ks7qDFpIaMINYxpPJx9Xkr
8lbxb9QQrm7iPb+ma8NzhuVyBRpAU+LpyUN3ugh4Dh8Ed64vz4kMjKo1XFLHuJxF4GB0WK0mu0l5
8eipi7BZ4Pznw1ZVP/Q5AixS82n5SnbNnFyK2c+0/REj5QSLG1dd8S93kCyO7mu8QEmZvXslhkRy
SKU4CC76aZHSVBqVbbY1pqXsHrPrjNEmk6o60p+XvINStFLOPt91wp2Ip/IuliJtQeCuxlyKHpw9
S/Xssj0sk3cd0EOFsZm3J5YCPRSr6NGFDRUeotU+R+elJ7hYSDl08d2vO4OBvcIuHHmTVeE0XcIf
8jHWMBpvSMYY7JgjcHKyklLGbeNZCkVfDBF2pfQ0bnvOxK0to1UlQN7Tbo7EKg+gd0mnlHreLMVy
CGeoCs71FULGCDm9LmQX9irzIKcKN5i1IBXcIIxlk59oIeZOt3ukJ6/+ntCOYryqpIToZdTuXXRV
/LZ0ThkuiqdhAauXLDuIE4UjzUmAWTRQ/iRHa/neDM7XZUahIVz1Cif2l8bc5NxJeSWPWet8Hnn7
vSqPTfpOmiIuMn4A9dTXg03C9OcB8J7eC1uZaWEWhORSG/T3K/3W7YsBFJ1HNhsubJQQixnrCx8Y
4iQojiQrHZlIHyUZta7J3ZSZjHebGRwMLGX8wKoKGFOub0q5AthGlLCE+d4/MMVq+53HxBdiuySN
roGD9uCwuDG8+M47Au7JNvQ2Gm0wOUHa2joGFtPXc9gmaTi2rXVZP6P30dFbDeMzM8eA21y3gIax
JGny7QDOzJWjImUmnyzAoqqnP8fbTWFA2uukfkDmRad/gl8l/bA7+YNwD46r/HWPMr6frXuktBY7
OmJGxoZqfmcx4V3wd2nWyW1vtKPrGLodJe8hxnZ9xstwds4tXPy44crNu1AtaIa0rV9jTVXttgCQ
iAgYQRRr+l8Q1Q8LEGdViek2zCI2ti39qMb9wDNBDVsw2M16ziC+1hTq+QmPCmKetVFk1iG9+tvG
UtkEEAc+lUAwM3ECeUN0RR3z31bdvRyucdwmscVTbUbcqNi8lxSDbanOWiIsC3SGcVQAr7PXz17e
AV19tu3qnT3aUf2qu6eZribFe7cA7e573rqN8FlOu8zKYhNuclSit2NfvwYlx8G97+fPW16Jiq5y
4E4Jq9DpbDxG9HZKMk+4HPfZGKIGt2w5GTiQw84sezWaq9MW2qfw4joGQ7HAQvJBb/QTIj/aBuTM
Z8uMqsnupNKWdX1U5EIve0AU2Inj3zsdR/+zbAjd/o5sSVUf8wbeM7mlmyjunpqxfJNzdSRcRRwp
Glzma4aQjGh+WOvZzvVQ5afkYzS3YPWcmtFVGTDbwEuSXJBqAjDdBjDiIs8fpWotc95hjXhH7yAH
Ekgtx1TJR5RFUoCb/MKVx1aBFTRZfm3uEoKlcKiGxirnRdG/MXEZD+7wpVFiRPqEGLeXyGFrfJaT
3ioM8gvs3kFV9nzpAfW4Z0CTErHMwLAiYdMCqL6TeZHH0ENXm7HeH2/Eu6BJHO0q5F/xxIYYzwJi
7DRlovl9dqw93n42MihRrd5n7xoFypuj1O0MJPKzp0H7oODZDszwpIh8wcLGgZXZzzCj8T363Ip+
/320bEn3OrdpVWAeYwTQBHvifFnFXfO2rNsj1s9rcDVitglWYkDI0PMs30zUamGf5Lb7Yd0Qjt4D
+YZbOGPr59glghQc1sLZl5YMJWdP/kd/onLYw0OnrM/Rekk1Z0zpxoodWlX8HH+lKvQjeY8IfGNo
o+BXB8w8L9up5W+bqsZdk9myRb6JCge/OlvpdUhyVZF246rT0h8JprGWLzLgxiER3LYdemIDt6G3
iE54cefKy8H+kCQm2Psdi3WJYjY1uSwmYAk6Z3ol1jxEMmpTs0YeGuE7HIfDhHbAgyyI3KpV1sDN
E31OZYpOPN838pZIQrdnACAVIPhtCGQ1T1ef0aDjgbZqLZFSeIIudbVw1lTsaS9zlIt2NqqMeurd
PN++YG5kYguMlWq34mmZ7qBXlJLw718/tYZaSm/5NW1UphWjis+LrDfhtcoov5OUo3oSHLZk6HZq
/DtO5pl+d8z0NiDgnV8XdV9DtkXQxqJKJbUPYyzsI7GpGnk3pj+9Ir/F3rD0dJuQGHClP0Wx5DpA
mPrAhTmq+gI0FAe/Ms6OALBIUYS7pf9Fc6bDlqdTSlmREeNiNMTBrxbT2fmYzXnSrAxQizm4L0R/
RT2XJaaVjsxK+eLxlvWu3v3/hp8dYo0v14Z3sqGH6t5GSPFKj2sESh9gY3A6VcXQ61BP5IJVaNyV
39FsfS5Sayx+lzWgt2NWPm4aRGt7cMvKscx9nMfh4yH4U6O/xjYzf/oWcI2AZndpHC0JVsT0qb9O
+B1gswCFX4j2krAF5QbluTKxkDEilqSwKq6IyGPvObbNkQqm/6+l6QfzfBjilf306brWA0avGiup
jiBIDSyBljYougbb/UFdvHeO9KDyg5ZsMUkHOzvSDGpbBv6wxyD19qhsQfvHifbTrkzXSeHBmnQR
T7LiQrHRG3k9XrA2o8AzhOByfzjqN7trYKNvzvw3npIF/WiiQyL1YwVJA9f6Rf8TJPp6bGXPBsD2
p/Ko5kde+DXiK1VfNXa2YTqKYH69Yd8j/RJouBY8ugKv1febfFF+DOya169gkuQm5O8IYvZ302dt
OwHrwbrAHNLb55zo8HpwSyjOgko0U6dT9DRz8F1gMs8v5ejbKPJGaJkkdI5cgZrfb1XyHmruRJz1
klyKGtqXbT6KHP8PZIEacXBPTk+x8WOnCVAEho/dqyxKiSI6U3Hn95FfqTOzsXigty/UFnLUgn65
yjFrRAe+jS7Tyjo3Cb+MpWfysMUSaCz1/atDZQyBMwHEoWXHsbtqIoRr8OJrqPMOYeCZoD9dzhwA
omx15l7conD4h2Z8ujikg22gb6k9ipsFhaj6bLMQJ2OutGRTJUrhgZYhC0zt/8IYuanZ5ULY//5Q
7tKCoNYeBrRY0o6A4T9pqcj8Ab2X2i3gDjBWoGdYtxasvGRINOUPcTZmyNr4979Cik+zyZCa4GvB
GZhYSYLvdqMMIaXNOKafGmAZLXWVFFUuYVsx1dMKFFQFBj9a2Qdf+tBTajKfKL4RSy3z0J1/hFxQ
FbcV5KhBkbS4jggWEjIgd/aaMPvwYBRiDUF94eVUNN3o94j5EzY/FOLCdOaJyeeER7d1g5vVO3Z+
RCrKuqzwI59/U1eJrwrWSVRxW2SIQ+aAVMNizUfM9Vk72qBYaAEsGfTa0Jq/oDS1YghUMJsm5q5S
AshB2FcC/Zjpen7sa8eDEq8wvcodFieUWFgBe1FZNoS/Mnab9OFT9VmD3vNDBxCLIkqSW6j7mdsv
MvU2jkNPHMfIlcVKGs75D4pqNl2IFgBQ8SVR5XLKjYiip2SVd4hkJOok5pWzY5T8I8hYWCejdOLC
mnOQ6gkbcgm7UXeCjwElTeWg5zMB81lmsPCoaIAmB7kVxIPNHfJNPudE+IsUrTDQsOVO74eoH0tR
H/N4CfVOmBL2+mwGWMBoWBtqdGUdJXKSQGJ6aQ/+7ajQZyATtKIE+8QSPD6Osx+PGwVeHN1yqYZE
vCNAnteyMNHHtFNFunyUw03XciH/c+wDpdKlTL0WZRB9dW/pzXCctKjotwZVG/mzvC9u1izZNKh6
h43alSgkES847Ot8B2vbi04EzoLH/nSqbPu7dZleiVycCvDl51FJMSuvMnx8n1KSTAIYGzvslVxv
aFPkKt9BYKXsiUqnvECKdMgU5kw+cRgW8RJGYcAvoeHhGk/tgvPz5wvw0X79Raq9SJPIuR5SEeeP
SY/ibojm/JqtoP5thN8BJGyUlep8ym/RtNbIqBL5pAzD9ofCg8JSvjyLW8+dzRHl5JKQVSSrWbGg
wV1+O+wqK4D1kD2jJ3KR10E/H3730VL8BeTSIKgqLf+J373RzD3s5/KwxW2+aXmVq14tHDpcuhqM
aWpMBWrqtB/7TWuG6PhRTY+fpCRWhJCkw2QO+Js/K4pWWE+4EBecPF23L86Kpwd09KRS4oFBJ4p5
SYDw0f8l6he4UQKSvMmYWI1e+xAv+ICpjLEUIvePBZfiFDaxC/5Acuv4El2dco2tLpbJGvueu9hz
5tPxw1NnsRwkm1Ugi0wqCcCyIudgWax2L5HPB6Va7q4GFibNuEfVDcdGiOIHrUbNadZVHZxaIU0s
/g2ZN9hgUwEyJ2xoftMBPp4bGH8pz4m2FAwp/xxJkljQ52D//XIkRfculP0FuaRZ/mmDujEDzTf8
Ruv9NZyCkOSXcD/oxIk5PX/30Vz3Vc2koCG+6hO47Vsk8qVJHmoRq0Ji61xPBS0zUhUfJq+N8aGb
1oqVkEicRaFoFfWKEmkei00HtGsTvNlUQ0E4m3o5pFRtaP/DwNf809d/iD1BvLm+/Uk9lOLvnKUr
34E9L+XWu2OTYonK29S0kJnhpUC4VEG4hHYYB5U7Ojl7c1/S9bVduyjGwor57yF615GrCycDts0N
vfeH4p2eOc9n7KJINtuq8CmggKWAgyc2K+8E4BDRZkzKdi2eOvLy3niDSge3vJaE2TK2hsajTu5A
KnlwQr17lRzryWZXOTNO0RzbTnbyLJBKRxZWMat+24clstFoM2FJKZsj3fOJ4UHf8FDBS4r+Bx4P
cwnclyWGMdY/5hcau9LKgF0jgi6kfGkPIVK8Dv5f4LTE1fV0oCIQtzcdwvHG+Ei51aT5h0K2DOv1
rXdPg2iAcO7/ftGJODikNvlmuvFAduYg1P7yI30HEaZOZgVRbp/MnygMBjfoh8DemzwudVlbuqbZ
MWVe/Bz+ppNh8qH+2cjAG1XUAbjmQ1kT/5Znc5il3XyTZz5BHwzLq2L2/AFX6CSYEPa3Q9OX+vB4
wELI5akxYp15AKDe5/IhwhYI4I0JOIv+22z5PjFaL1WxewubtEGO6IcXnYM7VttvKXEnKXQjMqv4
9LONavdT2pvOfcO/kJtbHWtWpQ0BANOUNzj/DRhpRKuk5Cs1GxdwddknxL1apkyc/hgWk+2cOf3/
XecxxH557d9XlSAqlaZcTkIRkLLEmLBi9aBDbEfGA+Al7AVeeDeQA3z1zQocG90VLX7vU4/HmkRA
s5BmD1ad56e03cNt0/s0LuNW/00kU6mK07LET0EfjtPD7SMpoRptbUnyMSyLbRdpw4/ejpkSFqV2
Qx+D1wLtpMLrKAJ8LzYp3eAKs5GeNHtfiaie3CyS6z5pCVHDQlAvFgeHECn8ROnbdNzvyGq2apgj
qqJMSNsKkp/sAC15SDrhQ+EUlT/bZ/3vpGur8IxZcKGaafcak07LIosH4Q5ZxlFrwBPGcmkZvC4A
2EGBBFh665DyEMWYN0zs/40Yb+68K3XIqSkwx0uSfrrynt4oYqB0upLDUnmeM17bywu3lxhUWnow
pRv3997Jd6g3lYZcG5l5xsVv5ESV06F4VChbZZrY1dj6ynW/7M48PTE57KOiQY9ywGCUD8HEL0BR
NuoDJPnVVBXQFiYNervN2BQVWbermigWT0e2nfFrhWMrHHE8NPMFBV32/hT91C54NTbGCS1LHTxo
fgFQ8oQWzvWlDCPqOT/vk0ZdOqB/HEZDb2Y5mRjJGDGpIwTQnu6Oxg5n7GO27f0V49On2U4NIPcI
YTxWZ3WpOsi6jgnhQ3EApE4JEz7YUHs3ISMRrGXNShzqT7BqiA6SW2lJCgjE+YjMvkijpxmGNGoN
OVbnBVetEZR9ogBJFu1xJ9Z+wDNAXgH1Lh67ONxUPw3SKR9qXUgKtlPx1y3nqZdHcWndTf15la3y
buBbsbVpdLckG6yz33iGCpbyPiWl7XqZW3DubeV6D5auwh/sSxF/kLJwmzrgr86iK3qkChsFWd6r
VCCz+FHgUFzFrgQTRl/FTz6GpRTJ9Md4MJISNuEjDMbZwbBXkmu33zLqbnLkzFV9jVIcLtbGKZPE
AZdrzoC3UPRnH/SfwlwjdXDIVsmxXDxO9FmF27mxVa4lcGqh72zM7gBCTJyi62ewdNxliDuSPlEa
eAr60ot3oYZD8VfeDNtCUt44V5smPe7RAAHCrCd8q06AMZmrTJ5jbo1qr6bQO2Cf1rPV1i51HKPI
RURQYJMTLKTbB76DkKjOxqc1Rkgei7ptFwQkN48jdJsQcgRBXpjjgCZEmcyO+5mRYqZT4i290hkY
HYTDMorR+9qhwGpzGulIdgI+fphr6d8vsEf9KZaJ7pwlR1rBkGdVa7HpYxcGB9xZsuy62OT4eGY7
NV+Vn3+gkNjOdNFsW3vJybvtRyh0cq4znZN35ZIkY3WJk8WDSPVavwuphqfIG/dRxN9JsPGsER1L
2jgvz5rJ+pKWagDqI15cE3dWiQfBZRtEm70uFyeRNYzQ6QeLRFXJHsZfJQLpTzzJZdrms2ObOLvs
m2MMs4tCWJg26uX/s/IJZMWKGankzRCbsD4WvpqLuOpKp34C6QZxijuMeiECjxGSVOPC6RcxT/SJ
FVCo2BdZUFgEHoVN43oZ7NkHTtqw6vgt9zbVlTJcxf8nv0S0Etw43+MYurBBfYTbbKXaX4JIdETf
+6GhUa3yxEgNeuVdNtuG+YbqiTCq9WdK/GydTydHMuL3MvBf5a47Rch+Oq2qgK3mulbmUzI+ZMOS
PsZQCECFn3YreyOkTVzFSYo0T2ALm4qtQTU2njU5e7tv+i8xDNyxSoyag8cRHudTLmxn/FQqHKpG
kMzbMT1dDuBRl6EZpkEVUmWDKQonPNKP/HkCIRFPXgKk3LnZqok8kilhU8xa/88THmNZp3/5tIn7
OChL+PuzcB6dWJiJEx3RctYorQb3bJmuBaPOT7bIFgx9NtCrwPyuw5SmUZuTKT98D+Gnkkt2jb/p
w4q2V2wRVl4xlJv0cGWNHYX+fWi5dMVQGP6RR1BF1ruc878b6Jhth1lqHk3jlhVu9EGZ+HqjouFh
yUnhZmCFKsJ6k/y/Uj9scA9+WdDR05/GYCFgAsmfzebendkGnUIC3IyYj0Ae3shfrM08NVCTVhya
enEjjYWbhTl44nrZbYmEHQ6pWdOgnNSY1kg1J7hbn1jvVal+GYMrbYy1uFnjOwWaZGvGxsFdMyvv
ERYGM6W2rwaAaa7QYDzz8Ftf4GkV56Bz33ZaAXQT6L7xFv/4wPpfbO0cCTzzbNCBWu+cfb5xR4QM
uTnDhi1nb80oN+TaZoKiVkMkl0fkbxvnXcPRhQpV0FA7PYQEV9AWSlgwbuMdwzOKuQ1YcRFIDiGY
qlrYYyt+TS9VWD/tcZ2/p8776Pm72yqkSV6FwG9vbZE0wJhyNRFhl5xx9OFP1qcmbHN/Sa/3SseK
t/dDajwbrAz4HZ6c2/14MmGa/kM+v5+lqaVAI55wU5dZEH7ry9pqzUrTsE81buv3320ChIWu1WrJ
FVGa/9DS7lsnljUSBepnUTArBo07pseMu2L91RzoLGms7k6Y3KDUIWcfozU1M90nMfAAR/YmmNTz
r79yhcm2J+31ccrMbVrQwhA/CXWEBweMsNvvDXMaMrqeg2/iI3AsJ+e0MefalJbZyFhV1//QM05z
0oNnRB7WZhHhk52u2EeuS6GHB7GdxNyDHQH/GQBPJ1CYq7M0+7c2RAtuE9p78mG1OLEYteSWONgE
mPk+RCb9tJjGQzohbsmPg0BZmrPsp4a/hEzVsuZGJEfshbUip/ppghLtrIv/Jp3rdGefKOmLat37
SQ2qtZ6RwtlA7oRj03ix/7bw5RIcWDJavXY9pmRkpe6IUCkgYshW8D9ABAX5h6YSJ9xsTZDH7byN
z0I7XQqCbBReXXHaxRr3hNNG8eh4/RPShLv9hKBjyPWCum3qpJfqqld4j4vaO1PV6vV89tjxQAlW
Rsz31l5tMX+FCKUeolo7Hr4MR28LwRZ3VlF+8Y6/8Q18GmOkNdYODyUr+X1DITqQNeui1DmiQzmo
pesoP7k6Uzyt5OvkqJB1OI9tBMO6X63MwjlhtHKQAwQKMrB+sSMQMZQEP3IRga7aFj/LPT8eCzDd
GYl7YL+lY8jM2Wi5RrDbSQKaiC60l3tGVOtb2SONmk/+PZI+ttUVEH+PXiy5qRZwQTa04Mvup0FF
z+nXm0yXPSiFVqdJO5WrwOHDosSbJhAzCMFIerkXVXXmWlhFPjqrpfTGjqyInkEkh7L5oW4uJ7m/
hInEmESWA22aX7EqDYF26kg8gJI8/tw1BKnuGr+XIbPXCFvX9PwMjGZgT5/CPBPMaRJB/tlWNBqI
oF4vGJ9qjW9ACkb4yRHldjjCo+qmafrs3UYblpKyZ5am5NbhMH8av4Gbup5JZTeoDs1NxU803pSc
sDKMAKFYw5SjmVnUX5DPp8MZsGmCaetAtF1Us7G5j/rcEElbAoQEthgyGu74zAu8eM+w0wWaovWE
3WSY/oy1++2Q2jbpc/E7pZgWq3fjO2LmPARiRUs3uNHo99M/CI46qwFb/qVSQRiCfzmxg4fz5vm0
JXLo0xazKQJLW7xehpeZgXXjHPQxVVr6Dj/ZY72/SXSan5jYwJrOjmwgI1jPkpnp9TMLOZT2TD8Q
RbXBT+i4DIL9Y9JieXRUmH0ySZSZldRb7tH4ncoDYZXhCiSk0Lave5Ff6LfLuJ4DPgt4HScTMvv3
2i9cows+Ti5mpkWIvErL6yypACoTs1fhQXcIgPbHSAQXtRTVEZJbSMIbsmxgLluXTNXr3HhSJHGr
iPYauInrpit/7+HuQqN+Yw8v4VWn607fDla/fGx2Du3yrs6YsMS4lhZcRghFeujWBtEqgpakLM+D
aw8i2QqD7JGZ6TYhAr9jxGFPxonaAExA8slBrU4smvDHMFJXDCCDdtxEoU+V4o24asTL8xE1/hPx
Ko5NIxP6lDxNoGVCl/2+iY4WOTu/n68yQN2b5buLW8pHIbB6NcNcZ2VBCYuCMZtrNhgfvdURG3YV
4vJZRAPS9X7tVLA6i2PAoneKOzl5uYbCC3R7m5ttGrD/dCnCPox9YAPbTKUTOXu47eyJRYbgUHBP
Re926Jcnz9lh9GcXMCYzKTNEe8BAVOvYlDplo2pSR17Fms2Pe/GcxRrBYjch8uXtEfQgz4KCicDx
cqLd3w7VuWaeOP58AeqN8z86Ol5tWZsoIids1oIbmjDRQRp2rNXCbnzembTSCDSJhxPTH+Tw3TZj
mI+upAjcpaGjWpeLfx633s7jlwdcyZsTE6OWtezFPlvtiKdp8oa1q4jPyMwPzgd11TMxRjIWhDMH
PVh04PwG1A/biwspFNPiF8pkeKlZnx5eOZM6S1RQAALE3D5TfoPkMO8A2RGVpTb+fPv7cLcT4Ubq
TjbGvfu/5fTWudNF+9nNOKB4jll2zs3puR99Rvzuara2L259BX2rYUJCdFQBdxYEZ8nBuFR+MPxn
Ckqns9WWKl/BVsdp/OenGj4LvHyXhiyfzMqTRM7oOrktpDiMcZYqHNv2+EQuXxELuAOQar4/akvL
FVjcOtWdANqlKGTVl4mnzd5CFq6QjeEn9q6CKfXOEMsUOnmadPWbpDD24MHX4p2rNZ4iy2AdJyNG
vIXLgV8WKwwacpKJrNP0BSx3VWAvunsz54G4xXuTPoeTELYDXeuuc0JcjUIqH+4Ug5L4iSeOe6z7
Amt30Fz9ZZcUke5JXie4l272UlbEUpNWDoKzDKP7BgiGcx6Wf7tVXE+K9KLPR8kaKbxgW5rNGBZM
aXb0hdTyBlQln+08nSrXD8nXtFYK3Jqp5iA5wVTWiYreeVOtgL09+ZOdl8evktHNJhGIgZ2QpwmY
d5np02vh4me1M0MAcRXoqGa46ylT0X0gswa5BlF/dgxB+3NZCQMYaCceteBVSie9kJiRopVl1SGk
2TQCzEstpDkA2JypCrTiHrbYcSG+EKvtih3/Ufs4r5+2InRkAoagf1Bqt4A4uez/YDxdWwX5NSo2
Na/LB80FhB0+gT3jxYvK2j6LDIT9dKKnWB4P2XPEjOQrSHmv9oDDuP4pxw8HWPJFrGnp0Ie+HQAO
w6y1AUa2PyjWHm8KDHlO+svrpse6YoIDsv4nMDvPiUPFhQOhNDCS5DR3T4751MNB4gStvzjr2+CV
nhM1NXuNSryJ2ilh1punv0HHp0DbZXet7qFHjLZgBqE3oAzhS1FA0KcmHLy3qC1nObsUVfmgCTGs
hU9e+O4r8zVPSzCMpF26EogHaeyokpPmTN6T79KckiGg7MRz0hvJ3ESgIeZXQN4WbBZQAZObbZb7
T92NI0dlg2zWGAIcrZ7QmyJMbNNG6t2iZad15pNKnjvzDrw2CibaeNlF1Smr56JdMFjY2Woe/O9U
Ge59a7w+TqdQCvbS+SVWwnsnIMkc2dhxSspi0EW8scaeiXMjGRLuQIFgjl7yBaDfwMgaukjidUkI
k9NvFQTXPL+Aq+9L1knNPeosBJNyTURTepuWNWOh+VUq7Vf5jeC7KidsOjuo/cA2xzVfcoS27q5w
KrRHri54dUbJLKkAcM6iPH//vilLlZg+RF3eHImx2uf0DR7Gl7diHFvrNpo4SS58PPrGhjTXPJLu
vfQnj9ejtFGJI6Kt0IaAZ0ik/CoPljogORTLz5bHqVfleWDSaAJyeLNPtVGIxun8qhlLl2UUuS1N
lU1ynBFiCvH2JW2pxT5k/OMc7rz0j/OXFJAp/wfK8Oair6Wq7vUJ9+e3K8sV/3Uq8OASg8WdANRS
ejO7hvFDobvfizeFvOHoOwvKk0/ERVGbIcMFMFj7NesbqjHA8+E+CazP/cUtAFKRcq8zuoIQb2Zz
dzJ+LT1q6cO5/v0PFnwHUOnOA39QtDXjd9Jsc8R8UV40ThXkxjPKFC7aD31KYlOXyqASMMqLTSbN
6VORLjv6i0MJNibcddIiB4CtWV/m7a64hvnmXVZpKN/To6lSw5Wz5ZFs+c4Cs/DRB5wDW7danEKH
MhgXgfH3qxfm9G+/+Wgmfcq95Q8NB/wAPYPDuCGa7UijYj8Z8F8GMbdqv8mzwZWrnJxeJE3lB/e5
bPQjiWYdZLNmsGYzhG7bLdsFmzbP1kr1brLQ3ZWkieJS1C1rQEg5fWkjj64GWkopzLZ5cqejFZ6J
izKhPoljOhYYZ191I1oamHlW3FbBgL4h/VBgncZ0YuwioCHiv78IMhdc+LfGm4n4uY+G/nTJA5DW
aeZKTpmxrg+/3PEc6CRCOBslca+DYSTNtr/ESRX+FkmePPlti6OqAi4ZONWB9aSvf4h7pRPmARKe
P9GGQar82Io56fWxIpNVAVRwdkPWfdwhsuZaQ6r5tMGOVcEyUGH6/ciyHLdDyDm+z/fHYrsqxvH+
Hdlp/E3ZdObNXP8EY1Zj9N5UDhpkLNzs6xtgExCHLq2/bVQQ4ew9oIUZMV6PJvM8tiwgOUoubcHw
yYaXf5nMdoqSP8e5zfsbEmW6I9bQDd1mszoN3FDt01g+TPc0t77XuoPLkeGBoxLJhZR2EuztqsOh
CkbTp7HscN/27kgXs7xE0fRMV6xRoydIoAApI8Guy/bPiXqnSCDHl8tEhr7GmsCc5AocyXG95lYU
MmchdEQFh+4tVmdTELy2qvk2BCTe4eokSwk+n8lbYdZaXYYBNtB81VNObWkC6sWTyxb9cM/UNnIM
wm3LEr9vtQ36NctUtOP1q85lRTT3TeWpWMvdFwQajcCNjnAm4AKGFerLewZE0gk358nKgobhYksb
yg1L+QAenvbI7fOanu9Yzv1oYSp2ayL1lE071KV3DRBHUXxAwURMBhqZDVayfeSu7sK/Mus/alQe
yZaWnzMMGEXX7N5RdM6hcGUs8zRJ+3V4x6+Tr8JSdgAm8M71a+6AOU5F6K3oRp5SdqSxE81Ko2vr
XcVzC8g6DYlx/zJx8lat/uRxxAYjsSLEZYKqQY9vr7UBEcurWrXlEVjn+YxC97jtV1I2Zm9WPhSb
B2YV+AAQAtOD4LP0rh4Ok9a7kslFsLblL8IF7O8SggIODReLPdTaZVEANwqRmNNhW6URj2oMUoJw
wFb4nOkzn9W8Z/0+ocS4xU3HkEpdDvd9LguxvoCEKKmkKnVgVZHtDab3a2rRPxhzToepZn9GzfiE
zx0auspMrzBDuTN57TLwNuRv9lURlssFxaR40CG6lVx5NqSMihH1+mSOH7m9+bTnPzG31go/ujtR
SC7oO5muRKZH0UYIUUsBzN3++AQ0SHkvyctdlQIw6WRejFbJVMfwqvLlavsKI+ajb7JEgzALC5Va
Sqy2i+Q/JPX7oI9F9SOUgTQ/qDuW5Jk62s5w241JzysOwSbR112b3TRqFpkL7uiBKR/NM/wvueEN
vA3mmfy6A/zQsjz91j/JEJFSL3GpLibaDWVLI+tf0mmaahJtUdqL5UsP12d/kOsJAO1SNqlwbfEc
l6y5JljcBCZzZWuDuf4k0ptaSf/FaDDjrAKT4NZZvq9eLxJKMG32erFaTF7Lhc6SyPz1OfOCnHYO
PlDtv34rzD7wKO6JvprrchRpihaX9l/j4aleVM8dSb2RqMEOoTi6TKdTsXO7aYnT/0eaxCgcZAQ7
aTI/5fjnjzXOoe1FyAL0JNt9CbfH4ahd8R7eB4ladUwMj2pZj0L00MiIdmbJD7rrFFkrQwtChTcr
OteBS+0ouSxpjF5+a7twE0AQpEXrPhwYhIO4UdCG2Vxe449X7etuAXfvPqqxfT/j1FPRFzJd/ted
uFbxZLIdtHwu3dLo8haR71CnxzfrvvhfydiKGoE/4SGLpJeDLXl1y7Fkii0+pyUFCL0FLkY6B7bS
mlGKpBIKV4zoCtBo30PgfwfDPwpduDpPkt9kpULSuuIkPh1lER7FTHIKgbo56XLLrrFZ6Bb3Rilg
QGCcegwF0Y+7XZGrLiagmaoWOsFWsU2rbm+zB3juSaBaF6cs9KFgd8dXZJDLuufwY5yR7ej+xPL6
wrR3o/TRYo2/PYBCbR0GMvsD10TgZb3bxwsAy06RoMy+gxMGjT7cv3Xtv2B8vSPkiAqP/en6mUgj
dDfJAWZMpdVEZD6HtT3ZioZCyKWLKxTlJWErsGrFrmegwrU3pRX4aOyBsbe7Lfg4MKxZZ1THE523
d++Cq4bzBevl39TOrja4JVC85I/r2duB66o2g+CHoKaQi/U2KbTjyPC4x42KNWL8Y3eMYSHPLJyI
HoWXi1oUQqHd8CJG5p3NY7HHPoPhhk00xwedKkiqqK+GgADfxW79JfRuDpBCrlYhbdUvqW/6rk5G
Y+jGy7iZ9urCUXigrJHCQiRi7ZpGK/UsYHDOlu0DeogGSX1+6VvhiGOXElbJIgiIGYNE+HsL9sFq
oU97g2cqCg7dDwUYNFyNNREIQOkKyh68Nagl5nuLDwytE7l4vWIgPNXeWxdp78eVXuNvcowWAZJl
eQZlGDJJEgUMxeL67GpqLV5kP5D8One9u+cgXWgS2WaLLloXg5Ryuwvs4hOyK0RpIdrvdgoNw/QF
R9wEt7LUGUv9aj+nm17pVKuotJHJNrqfr1V2esMYav6mwGjBMTZj3A2KXMWJGQb4VsLBUbsDpHoP
YiRcHnOS7KZNPF642NI8Gtq++b9cXCdaKqvyETXquYUQp8BgjK2ptMWDwP0qyyKdtbjDSYvdfdXF
SmiiAhkXzDoN9JXTgXd0gOWDskAeGOS60K5W6SbPAACjiLOpD3lOsLBvlE+Bu/+8nXqRlcL1PPfd
HuXqDOZJywMYRSm7iJVdqKkYznr5XUyicHebayKK36B1CBIVOTwht8hfCdKaEAT1ttT3Dq8X3zN4
8YaGel2cukfEhd6E9sY/aqV33L8ftRjpb7JcqmG+kt1DRoQsXjYgXqFAYFlq83/Op19cZMGzgV9e
UnJZ1LNubQUvLD5aywlZumgJTUDfFxUzBgYY5e3x55g+GGJntSPbaILbDCBIrzdmigdiZ8vHdLFj
e8roCVLUJyZwasbihkfnEOxHgmlBrAT6J8HcadYJk5DNQGNGtzEQQXHVR9HSOXSPWWYbype3IIgX
EdH7jOBneY0extT2PHm0nTUIrpoCmdLFpB9NETItP/PWGUpjSWrUg1WkKjScGeUbWmhrvKxUf/Ts
Ws1TTH30H4gP/oiLQigt65y0SLX0vph334FM3Han7xlfjuZUVjezgghFgruCQfzG27uqRlTvgT6z
rSg4wV9ANKxwF/0nwe8RJVy8MYHjsjZRGpqGp2pPCwHdOulUTgtNbtEQEQ5F+bd8anzfpPpeIjia
cEjPlR40/T9x21sNYY4ZhsWsb+6KUOTUpGNkldUTUl1mOM33NSlR8AElZltrFbloA90spW0S2Abx
KE5ORl3s2Ws+KPeZRVvCQHZvW2O5TmgJv+yx6lawaOj1ZJ/QF65vBokjhNisI0vEgnTSVpofJ2HA
nBxhX7els1h++yQMy2qp6dJz4AkEitJAatY7zTKV/JsjQ2qS9dbNS9gq14FnX94dfZgpxtB3D1BP
bQPtJhw5zkfkNQz/JBLb/exRJ5N+GlcoMue9/W7xQc93aGToV3acUjwZKGwdFwi2Pr8Xwf3ENmP3
sqP0FAmLS9aE7AFNW3RJ5H/AFRSog3W0VeamgaKOKLLcapU19cUHeYhKdOjJOyxoqGx4jDMzbeJ+
Myg7X0sdt4XbEAGM0C78usRIwvpfNn+fMWflT817wpG3v1FuLKLQPjgIyEJO8naT1wzdgubwrXPQ
EzXiwB7ld1XOiCiEjYrM85B4bMedc4TYNtzBJ/hqp02plqJSNjCtEntO3OZkBC0p6oCyQmq81DLg
M1+tZxQrOdv/BQQmLOJ6LUVdzvKDjuq3B4DbHEuQT0hOUM1BlNzua9DClXNsuktjtK249+G21qjI
VCE1BQJTTE/XSrxobUmJ9CsOSNJNxPUyolx1UADorxxEeEHtFGokM7ySTCQ3VEnDtK7Pw2N/Y0X8
z1VpXDjeOFFWjh+V7389r8SdmzbBvC5IYJZe16e5xXjwSH0Xo6YLfZzh6nq698TGeh6FHgpD/v5d
A8xRUx7B5R8+jpSc3YdSTqfEh9a+Dw7GVbaDqmPGMxuFt054PPmt0kV2pw4q7CE980QFNkEQfN4v
I1bPl4nTBHiRAxjPsTwTtf99INuw+MmTDI9KqGvo2/JvcgwZn/q4Wyy/o/3lGZ7E1k/ll2RRB/ZE
iGWShIi2w4Kmzoez1VbK1uW2MNGQAA69jwJvkavPviQyjgqX9/vU31oEBqESyumtf90SBhfHOlM8
Tb8IjZi8+TxNCTDOscxlkphWtBFydsy+Uk+oAJOpbOBV4yXQqAJAoKpZ3r/Ds1r7ycMXRpVQxpZm
uuJfTFqriRGZekb7TWMZFtpF7qWuL61HDBKFKHda4sW9S+tZR7NIXtclXmbkPAbjjEFRpGrDO1Tm
FBPujQ7pbo1X7Vd+v3p+tOc4/48zYuhSKUtm7PWcds5o0X7xgGyA7U/aD2PJVSIg/H8l8rDQf21E
NVYyBd+wBznU9xpH71DWa4vPnWgh/lDy5P+MTDrD/6A4G/+pvFkWOISfAq9HdKXH3Bf9ZUoJCon5
IztN/o5t2q5NP81CBJWGln/z2lT5ygO0ZucY12ScDQJaBhqpBblMxMR3KMDyeJqw1GRBh5QmzQ9U
qIT6+d1e0QXxZ/SGPLeS3XkrThuZyd5PH4Fqh9KmY3S66AwPqAELveAZQSKjbK7kbXV+l69erSw2
gmBldh10hT9RnZrg31fnqkJDfB/cCepHobR+458q4JXbpPJQqxScEbhn39LBSGoghb3uccSGDtCZ
xeQZKLMGe/4rlxokeVFvy+ntExvK5XLWsekpxq6t5f+92fOJxNCanjKgLPNEiH0RvxgKEIEwAtzK
G4n/+YINQDBvVNlbPhtRqAglVYYbVzEreEcosFe8cIFduS7F2tk4aWWbYkHPObV7IywT9UxlEtAU
wXcdTC6hI6HM7doOXyaAN/rBZTiluq7TxQRKeEtVhxGuEYFJjYVerW23s2LDzI2SCbFbeJ2AmWsx
0bFUfU2TogpvzSHsDDoEEuX4Ht47a6x2j+SL813PpaipnFlSe70gomYJmLCZ2roRNJrF9Pg51UrY
UxLRkw10j8N8uPOHTs0rwKTPEupCQOsBXpwp/vIlMWDeyE9YDoCunq97QdXIbg+s2yRC7AhaSAWN
K4q4zF8rDC/jEAYqcSCXB+m0eGsZ5dNV0yZyfDbhLVJz0GHEoRj4fgPDsRET5eGi1JmGqBPV735Q
KPS7UOsvlDFyKc8boCjsc7bHYP/irrMO73duevsZmZB3oL6dFUVVPMMgo3x+MAVn14xqk5EM3W6e
LoSytLrRvbuaLO+eTTJc+IWkHTY4HLi1ORYz6eMBD77H6vxpWLNxSySMvP67eif4szFGWJ/6m29S
XonYZrBFGCdxpwoHZ/0ZIQk64GpphZnVxbbcFrmHdIcuJjddijnUz7mcR3grImdJGlBYAuuhQnaI
K6NCrA0uKF5OPh7grucWkXkc+eCgpIVVeN79d4R36jk+l3LFVr3QWr7yXp/+IRCFk6glXWF9VZ4q
IxQOgjYkU03WVO3Dm6/FLMOByEp9YOXt4HibEseXm7PZ+M8StnqP7/Lij5ZkP6I3iCRIEpazr/i5
lE4cc/R48lInjez3+Jpbh9b+NXDhgvRfex7Qjxr0DR4CrNdwSLTCPS9pSCHqYUuA+sKBt2TVyabo
3bs/D6dtlGF5uV8dMIsJxZ263e9oXtmrb2oPKVYYxOwgaFHOkrJxlPnCghgC/SxZ85uLDOSsY6gJ
TW8k9+PKzjWXH11k9Fjd95dv9FEy4d0b2TiYgwZuA8lAnNg+D7NV1geJCZgZ25g12/fkEHktvHSu
bBWWSfCqWGVjkgjE1H0l1viiMeAyTrAEru4pQDkzNE6AiKd0yUDjyuoDQ0mCpTyk9enz4l8YIS61
iynUMParismaMRnVHxxvGUrozMH6eK/hE4+5CvPhlS+9Y2p40kSQF+22gsD4yITRgFvZM/4/jka2
taamMoONigYTSHFVoe2u6yVo+cHSOQRoKLMRIiON0o+MXe+mK90j7UwIko5LelsVewxs8XHsCxrS
ze8No+d1v2gxORiJGBZBcF7K+Z6tZZCpvSyRL+FJMYbl1Uwsyb8e8zyI3Vu1UPKOD2CVI4tG3+Xo
UsSUjqMbO5MCRIp2Uu+bV2UBBfnsx4dxLIWGOFwifr7DWY5tf+E3teK5MaAy8xJJSTFSz3O9rISh
moo98+TOUNPdYKHdtGrGDbIq8ofJeUz82OMexdlZiQybd0ayI9i7i8XCx28VAHb0GI85WLarnjtP
x8Nq0I6XIDX/EuPjn/vE3FB3iZmruUBZR/+OFO9Y5loLZha/JaMC8Ryay2GJFDrTTpfCgk8zsr4z
8SMGsGL7AaRBo7dIR32Xvc4osY7XTxCmHXdUKfZ1B/KvAPquzFvTVuiBHjT3ADQD75BPnNLGDXpL
so1myT20D/hnmOTItNMw2nE1wQkhSNiSw3UoqaKFm99e/W+CbLqMBVDArcSRXF1488bklgBJYkqJ
SNfBrgCHDen0jH/w8hzlt2qic4P8LP+s5wsxHNECkMIcf9OY4Oy9prxM8K3hvLPs3Wik5pOEmDK/
SBn8nDCvVHyggty7WUiqEKOVnX5mkrfj5q4ZmJaDcigK+UPql+iVh1lFpVQRHZnQ2ngFpL+tIv4q
1CfdDqFqmYaw862kSX450atS/oi4GU5/poIpKriPGDQTpdgXNYQtakuL5ImVuTL2qoZFXF94ygkL
3KP0/3OO3Wcinmo6ISoAUjopEDcE6tZDePKIW7VH/9wWwOOG05W1PYzc/Rlfo+tQ2b9nFt1fFyNG
e1wkHTle4p2qgw1PhaNM2ucK8dxHrGc6nAJdOfwIUo+fmIuNEChGev4ixx2ruXcpvKuKDiV9qJrz
e2y3MeLoIQNf26kKOleNjhw7AivwhwkTOwOJW/yi6m/3f6NnFQVdlJsvlKaFTPhBglrBr+oahZKA
DXj0N2p8Ze8ntODFR2/eE3vzawoqND7DO+2AjvExT2XNf+ooOMFGgeA3d5PZC31TouvSNi1+wz9o
XQxIUc4WMHQy9sg6d5xYGgJG+fF3AEjs8RjIlxtlUpw5VAvx3WoldZ9GUWWOZu4qQd9i7JjzFpX6
bq8EEYHK3y78GeqzQ4YRUZ/D++vn9YfODJvOmZu1i6xjI+Ji8E/QsWNj+kRwAzHnxIKrzhR1lgch
Vqm+MLdS85LUnrnt87zmXTVn+8Ygy1wB1hD6I9i287cBmJtudHwy3xHfS96E6yS8jHQQNh/lEoyQ
MKb450WAf1nHTi4RjPxf3LOTJNJbvLbT6HdOWzfJuhW/lLG/PRprM7E4YIiIDRBb9RN9f/BydjWB
V+W+kNLBm5oASXF/uelBaUKenf+loJyzMKZYe2t5pPCNYcuY7aNfo3VNb6E7yuXBqk48dDmlJvYj
iGcQLR2wCXE2cf5N+1YeJ8fpV2BWU5SmAP7MbI+wZFyL4y8Vxmx9y6ZwpqO/jQ1bc5IldihNNKuy
15jF1zzjNc+QqBmaz9gKZRriLmF8XTsdcoyUvra4IqeDhr56nYZ2SK6JseDUjoQGDDuDROEkSarR
pVyiGqviW/aM5WUVT6gtYey7G52yQCnz0bbGJef79gPfMkNa8cdYdoQ9uOz5H1G4iNRs0+wZSmNe
4Vqr86YCg7jmK5eFDcRhDuzIZLnYoPHnsRS/y4vi8VpNcI4labDExaNe8nX8usSZu3kKuRV/5QEG
BTVF5Es+BO2QYH/iawqJOSwYzFgXMVRVddGWWG9sVr+gxEXfR4kX8f9hb+9UaUJCzoWQy0v24VCb
C8fmel52H9M9fVzcM0xJ1Ldbz142VWIMG8AT0CNx8Vv5vyTPP2kssIQqql0VyeeP/72ugtj0aLdY
Qr8sX86Y6N93jXGbZSegXVy2Xzm7JJX9+sP+GgsZ2em/QLQyhZE08s+V4xvaxlm3sTtFCU6D2k8B
DMFm3YZ1DcrjbYooglwnEPT/PD4/sTQh/LWvlXZTxu21UCYavNH+DbZUHt+z7OSm+ukdWhADcUQc
8suwzjfWIDnSdzu/OclhH/e6qozlbJY4KONpBU3eVbrxK2pRvVRnMCTTdgswJNemSFN5uPs7ERvQ
KQQf8t1cAMchpbZWp6t5rRRILBv8eP82aT+eRGiwyQVjtMaaWkAfpeosSxzUgJM/49nlot2AjGWh
uTJdPqDm4TSRWyfxg6zTillMKXV5TsHovP/x25MVVKkNPs7CT66jPxKtvqCq/q+ChzZUgnU4s/dT
f68IxAtWTFLgNfYgAT/pfAai+iW0G9cesO9DOtRcHAVGVrhwtcX6JdaNbUWWxnIN4kYGknqgBOva
Dy4XHS3VH//+9ojP13r0chUHOLN07DAoP6UjJGOoGiwbRudygCGyzJmLbIjBYoZukVvto0z36KXx
Kg6iTxbdClL1d5aHY6sjZN8g+swLNw3vaT19382YSzATCsccuQIm+Zu1ddU6/N9F2JQRPczzJV1g
+2jTJPvS/TwWVOIGMM6F0OwrynA0XAcAvDHLDUaHofb2JN3FLWOuQEN+lrwOgbbKrV77hGT8GuUz
gLm1NpFXgE5oLEdVsH9yWDy+dP6ire4+9idFabQJb1Wyw/WZMm4yl/QzwXwQoODrkIxqVMAqzww7
NbEGqCNSGkby6zOXddSy+bzV4jAnt7+UYSzpoa3nCPsGJBh3GKJQJVL54WDxZuuMFpuLIIbDTUip
wV2Lj6+FK2YgPqvSUihhJdqnyXbs5520lIks5uXMS97aXcvXNMR3k89XT4k+LBfrHAmtly4C/arz
C0kiNaCVqrWOHzrGXD3dZCqU0YiscZCqkWmn6Nv5jALDhgP7P174S9djksuKxC/FM6YRqedrA3wh
xr2EUOZqOd9kb1px9QSrkjCogekTIZhajA4gCKoOHlYgQK1NHHAm9nzh6l96Av1pWlG+VjYdP33I
IgAEMqGDN+s8vkVeRCkQ6eQRPbRomXzvJzucnETBz/M1ic7Wz6yJNHaYrC8nBuLn2vs5iOhxQ0UD
UhD43uYHAiavpDNvxkaeMdm5k6MDaNqf51T+Ic8nrwzyR3bZwNCIHbMHDMMOPl86fC+bPK3QvId/
XbEV+QVcXynX0jtc7MFuKiHx1u4q+HF80bLYR22+PD1JmGhEN969Eu9yyOwyzw7lVuu6GvfKqLFz
KU6Lw9SSLTC7N6fNh90c/dzFL28vlVxZOe7FfzZzKlL8belOMuyZPzr9Oc2a0SvEuySfLq9h7acP
Do7ujiGQdaKtgnwI/OiTukUGMzQal86c5Gs8IplrD93Q5Ng3aGZ74knk/0ETKn/+7B+Q161lQl9s
Kde5kSLilS4lkd3FdHAlPR0JkC65u9kTPGKq9gk0lbAD4cfYa3dZBUnYWTLKoVysmOTv0WXujU26
203XXgZjekQ8V5X0dPrxWlRUvx5Y2wIEnVOM8FVSKOVvIAeY3R1bYfdKJar5R3Iyv7iRLT+jaM4v
MSpKrOEQxK7RtHh+Owyb6rfuMC3RPY19lJmvS4ygCY6GtJ5hYt4eRzPtOF0tUQenuL/cpHCPLc7e
XihLJTKBYLkE59skAf6KFCUr5HRPGm6gqzsxMR+OSq4gCxf+7pLKnq/T75eaA38XNNSpUgCry7NL
8tShhGPdNy3GZBdQ3wNQCbFPyfR+NQ4Kl8dxYqcjz7HCyNPI/UCR1WnCPl5pk7qiYOu/UtvqS32K
sIXQ21FNWnDJFdW4DdMCM5gOYRgjeZMBMzf6tUORM4AuIx7MgCuAg74lI+KLBBnirWd5+vZeYC7K
D0cnn+0H+0WRDFO7mvzpxuHumfSqH0/cOW+QocT098UJwyPhO5S8yO9ZFdXiYj17sKxDAK4+jOK3
cxv5KrY2jnJ4CHzn6oZbv7BAuCfhAscvKZPIusL86TF1g2RSwWdi0mql/aKeiPhd5vFrCJSRx2eS
nypd6Dmj1xl4ClDnwC3aueK2TlC4aWIuZD4U7HKaFUoMVDxE4RbQAMvdi9d3npStx7m9PP6eMuub
jEpZndh2/RXe8vRrqPYuThWjL4SLS46SlkOPpSsRJSrqGFNdZDImQppLH4yP+BA9H0ibJGW+Uemn
Z/E/nWySfH/Cr+HHeY1H7LL9RfrM+5u4AgXlKtFcGaitYri/yX8p4UGyGjSVxcs2ucPf0ycrQZJ7
XKC/PaTsxfviUnpJGU39WNR5I22OXof0MXnVHHwguVrZC10K3xF7IPi7zWbtT2uexQA3VEOtVr+6
P/S0+cS5m9pwne21OKqzpSkEQOqs6uFB+1J9/ETUZo2m+xF1WLkk/qIP//eL1GI4kAhCfcx6Do6K
Ehg6V0Hn+rZXRqb8DgOGVJfXDoV6W1Kfq2wLPP5RRoDYif0RwD3Qqh3DQWc9vN2MEgleyaizcwY5
K+/yhtexc7t9wKc4ub0LNk11DrEkI4+Oi0l7lsAlbIjkvM5/flKMcbIdqmrGWA1k+ehgVwhudHNs
b2fupm9FulC/C12525AIs27hS+5SWzJEEL+n5K2wfwbC6msidtlR7JVipAmymZ1MVxkv84JdRnsA
AFNRKojb5JqIjQYFyIaqxAfqz/GneaDA/KL4rzgLSkjHG6dXCGOvbxyr1eIjnLIOSQ8Z+zEJfvxs
fKmvtjEk/ZuAM+yvrPS6t1zCmHD8HIqtvk6s1U5jog+RetQv38KE2fnVKbTirRQqE/SxdMZzxA32
Kp9s8qMep46EUSlRiksmBMX+iDWbvjP+HhNeptTr2ipR93d/VJ6Ebii5ARjZtr8/O10RZ+C3nCuK
v910e8cJUXyQbFFELcDb2agy4oekEab5h5AFgFEAPXJXlR+MhE7d+iLwj5+1TvG+lpdXBzotIurC
im01GKtXErXAX5IAYyyrK15Ko698Rc41mrFlvp0b5qhT/A7azmrJyB3jRuOBOuKqIECLX3hf79sS
4xVxCVMCY/DRDoz01OsVw7hqSnNudEBVur4PKKrazOn7ScHOJb7wN7XSz+PE5gTFs53OE3JVxfMr
fhzWwE0xNcb03vItqTRCm1P4Ez8HETK7G632Ubtj33g5uYsky245q4tNkCZsm1xuc1VJZqpyZgWe
WjlB8dMuet52dTkwZD77jTjlKygrNu/iXYPTgoqQIXV+y5aOW2NVKcF0GS/HxXMDmRO/QoxoZucb
GdpRrM9ZLRQwiGx3wW0cYX2h+vQFPIhqCvaUXN5u9J4E7whl7yPH+sZ5jkcDr6OkUTl8nhcQOjxr
zdIFDdwix+ZAmPGl3blusM6rdHWVCdQQFw6aMjnSXIqJxmQhr+RBtyirRd+V6SAUyR+IwXxOKWwg
SlnvT0v/yb2pK3BzAOMVyQztoqIjUC6s8e7jsLslZrQ3rT01kPljH0vpLS2HuOw03jTtf48KPpLT
Ow0kkyIWX4Me6sT7GbWbb57J323i4u21s4krPp7OOnE8n3LLEgbfqNHNLBaQf8Q+Xb3x8JKcMgqN
g7b7aSKo2unrxZRUTP65FEEv301vXAoiK9bHtYvkf3ma3iVjQVDmWmdXk2tKis2wPCCsJzapIOeB
tXj5IB++9mLHLNF0nwDy/Ogiu8+ggPTADwKInl35D15C/57REZS5kRFCOp+nAT8pYxhcTUoSU95X
unJS7lgfcX6uOfApLIyKdEyDEJ54jsd+iazRFHaB0G2Yt+QVBy/gpmHTWvUHQd8WKP3h5w/VHUQa
MH0pRE9VfN8UgX/0UXNfZaAF/f4SGl7frScXc/dhKz7kskcKl8FOUm/GFdgN/YMYLGQreJXN8JjD
8GBFW5DA3cJZd42GsJKD72pebUbmZquD/DVDZg7Ce0544E83fEd63mFd5dlEHf1p4y8+Yo2Lmdy6
LEu1aYKv0np48aURsu1e6DgeGlitaPBqy2TlYO1PpuUxW8tlMtfUvgs7oOUdbFRDFPWJbzTwx2zH
/72m6MPuVphbYiJILsuMuVaMPWqcoMgzkwBlenuVgoA5kYimBoBe+BJnzker9XcP09ZCv0li3b6+
TnQFoSDh0YknnyrLorQ5FM0TLMMPF7o6mBsXLd0HHr2lYiU7djK8XUEAsyt7Rw9ztacLJ6D+uXT0
1dTpkvKt4uggfURoZnFQGWyKpxL0/N4T6/psJOJtR7BvDoGOHywoN9DP6m0nfDS7z8gC5XVuBi63
PmGFdU3MtkuoBU+PXEx2xnlWX4hYBTs1SXrU//OuAzUi1NecxVoBo+F2dSMUdr3mwol0s+Nw3xPF
p9yYasufJFgXOjkNrPx1ltJfkB/nfyoknfAHvnkSAYeVppucsfELuY/W2rtl8K6bT7LtdfLjo0z9
JEvdkX3B2nUe7S+ItA0Vy8bC4Lf289QQL+XoJXmM2RSbeSJ7SBUtUXS/OIhwo5rCIzXcoAI+yzS9
xNvPc1rqa16DCgiQnQnVbMuh5oJ9N++q+MF52C8zTRhab0SwqggdHiRwONXhQdwR+KATi+vWR84L
RnSX1Y7TAeoZs0w0kaTkB2bPjUSKVcRsGMtGUcAecZMP+oXVhWcFvR/7ChNFyYkc6+EKo0cE8Prg
DNw1iedbb05MdxT9pdy2nTcVZ2k88XSrNIxF+uNRcwhTqEEiXE5ztzyu2hTwq0O6ebU3nU7hwIiB
ZaW1Yco9CyP1l88l5S6BD1TBZH92z6lFs/Os7X2u4VhOMIXPK845zHEF9mB6RjgDfeDxU0TAo9bn
SRbphisBpiiS/7Ui5vfjZGSQND7YSVro9PaQ//ucu0bsxwf7VHEJoMgplAqWravPiD3YbiOl7R93
S9jV5Icj5DbpsoB3DkmN6irDWlOTTtlhzSYQ0kWdeApiOXj8imoBLHPJrvIkH3ihYYI3QmHj8FE8
64RRFjAhEkRy8i+6oWk+kcPq7kYzpIFvEwk37RDGJnNrBGFlJQyp5wg+ykgzQw4YUwRuAokP0SK2
5rk6TH9djfUrobdZHp/yqHIcGawdArSWl9uN4dJ6W1o98af2F0/pv8ga6GxAODSG8nL9PpuHjfwI
SzAT2SbrNfuNeV3ntntaxs2cWKAXP81aOeOCWU36tSCo0BNuiNMMXRh/7Ek5F/C/uLydRvAEieOj
R1xqmphYxtpNVVL1u5oNU4h3v6iaiJynPOW8iwYp6qZ/zVRZi+lnxFidA1yD6bibKNK9xbgc8KuG
BetWWCdonWyICes4367HqBFz/0pK80dokApNofRCOoahA0tT8SojeFbKVwSPAvnwjvPx9xv1su3c
52vTlSGfckIf9cktXHSNm+ukPYb6aFm2dKAS/3eOEG/Tnnw00ShUhDGMTiBAkCwukmLRUWWGdPhC
9XhN64s+QPZFanTbcwfzasOFuV4AGHLoDXLh4WGkmwlbsLsxFLO1zQUZIuZyXsajkpEhY5gNxd4r
A2r7LXkmQ6nWi5SWQTVt5gyFHAS0SiYp1luteM8seRzcfUjzixiTQku6sf0f6QwNa3um2ot6T2lN
Afz08M5NLtx7HsKyQZbrRkwhTz9omCDp0Un5GSmBsrEVROjNuIx0lb94a+Cft9IjEgqD+KaIIYpz
ZoLKeU+Tao0Ui2CxPWKanELFJO1Owbqutms3SO95uXT3AClfJGWREBhqNE77slsN9F45lcDDRThv
7F0djG3rwjO/p8YKVjRs8n4HnDcQZZETzeEJ+ZH+YPVzsqvGO0DcFIRYiQEpjV7UpK8zgMaLv8I6
RWjPmbMbrFUs44yJA3ossOBfAN+4ucPHnnFg9ES8uNCk+cXysfg0ahaajuF11TmbTx+Iz6ArT8s1
4Gcjvw+3Axax96azW1i8p+C86K2RIEbfZ0Y/BysSCs1gRGAIYxWKIxrqjy41oDME6y+DMrQcnWxB
kfC8XfXTRMjtajxe5/cUo6eEWIXDh6RZG2U0mlRfv2D0IJxdB+mjKJgn28IooGVfLQ7vpzLO+miw
gJbeMqdZ2mHwFAcB6ej4eAeBL7Qfzti0sRJNFcArpD5LhXoPn7oYZKA3kmvziCqN8Xp6gc0yUgOo
7LpertsSa3IviLQoKaAhnSH2L56p4GbLcoKcD9NLZWJ+fZxWbmtAHZ7C/89DKeebX455b7h3L8Sm
Xgqi8oapXoIsPw+QdtMLjwPV01z9cKxNjFgV185TtjEZWeJvrwDPGS3kvnenK36Rz/W4HxpSPwUK
0sJhaZxzuHeFxlsy5YS20w1ZlwvR/CLCBAPVwiVKskgeGc2ijlzUlK8F5UJUCE2QuwTJMC3jbG36
Jliu1TSZnUyZW26kArpphpJ+0mLz72EONVdurbiM185s8CMyqvKofQnvq2Wl4Ilw72IIi5HObckR
Xp5xcIT98ygFTK8Myz9Ftd7s+Ix8g8kxxHPoRg0u2DvwHRJKjRzxJWqK5SEcfi2E/17ePud/sTCB
CJMUWYtUoGvoF2qWd+ajOl/9dNFKQM2pO2Hbmu5DGulO4dxKOaHRAz+R7hlOoarOGG3Ed012q7Cd
3oySigfz+QRlrJS/CGVSWUXmgkq/2Kdi+vYViqcUxMbRSDNtdwelN705Y+zbJxTMGw3bMw4T5e/Y
qzhZ2+OY4LW63SatkAPclbeUWHZ1nK9fbnjxE02YzJerEduMX4Dx50VcUzCwzg9lNZJbvCBYwD+5
8EuHBKEabGMuhth0qLCrKjdFZz6Vlf3o1fUdOaeDGQR0u5UuBaJbCYKsCvNjSzH0QON4S9qULSJr
v5ZRjWs3yhX2iSHsDopd2prjH98sZsyGzCdHFm6FN+lqTek+G4pzgeckvgV8fsvvGOLaP3+423XX
Q+mTP4PxeeWCyxndYjcEfLs7YXcrq1thcne38HQCRciTJVoGFzW0cPnz6aAs1TlLeX0Zc9EOxAGr
pVC4Lj+31fmXYO6SpLZ/kuTYR471mjkDvIpVW+TzS3zCt0w1Y8iNzjAOG+PYRO71fckki14rROU1
0oXqiS9SdtXBYiaeHwB6jNf0ICG46EjAKALqe67RlALjgcBHC5ZplMOlT/zgFchajgESdKrWR5go
H06wv2Dns+ib9WS+rgm2eqtJbChrJhf+IMHCdWaxrjcwFVH/CeeM9l4dZXudWTFT2ZQ/CKDBc5ri
nW7qP7lQTPCJF7dkwzkoUCycEyYViw9KzFkolzCwIRdvQ7HRJEBSPm8O0Cs8blu5LWG1mP6gHfmf
69OjYHx4pPNv7bRjlKzlMYh+dxvch6DY+S/ZhnoaGhA3FDpBDUN8/ifgGBt9jvdbmtK8+JgmadMX
z7MrLhYKYSdBXfxDIVonnCYhZm55adZH9aVcpiqMe8xtXGZ0RuMt5d24X95PmDcAVEYA59ZXtSRC
7/fWenINQHYsrRrFo7iAyYTHY4YznNu674Y/a8p1wfxvofYOl7bxoOunxEgvSrJys/m8lNwbGUc9
4/LwgvUfJsYyos2R+sUPA9C9UBEL041t99az3kUhA+7szeEeAvPR8rMQxGqYI5uW+O/orYFR0be2
izLTMdemG+A3x0azsKxXZllzKIX1OPKloBzlhjSs9iphGU71tLVBh1sZ061lvfQRK594DKMPktYH
OF1gZj/U9tXks2PW+6s3n3kI/5MqQLkDwACx6caIjvAQxetSb0VEKAeGbgT2m4E3lb+zVdlhDNzE
fYt+T1FzSCHbXdhUQrZ4RGiTO45/MvUt8BwPAiSscDhP4eBN7OaqphhH4KuLv3ieYTT2tfEtgWaW
RRaKuZWzjaAelgP08Mk0dpJ1DlUJEJonmbaFx0dEu28GXQofUCMuZJf9GzzQa+SxkJn07K1zHddO
qNA3HW2D4WtJYYH+dWMi8/oEBfTekqrHFwvOlYPyzS7PKfr+x6gmDbWbQH5/AqWqo9jgSC2O0xft
bseGm/IUEbQ75EVKnAgKoV+t9vP31kvvIr9Tc1TiVfc56u1ZbJgwNTaFFJZihMB0W390i6ZYkqy4
OrSWHAuXm3SLmHrpL+nRIDVf4yPomwkVQLJkS4vcfXFGh4fdCsmjO2+VITBOARLtghbtZpzTwNhT
zExYDXqqp0f5fiQkm+b65gI04fFo70hLrN5MZtCh8vyDy3Gav5IGVEB50e/3ZNONZbbs5FOSlCu6
hroAH5OZuRMMBXDsUnlq0O7CVUBozuZLeHkWIINvZUhWo8lZVmGr1l2vP08GleY6nlgMsn3L8S6c
zbN1wX3/5VPu/Z2MI9dXj9NuS8c9lvAoFRR5XTLlfXEYJpW5H8PmqCaPAYFnQrXAQzp5kRyP4Fyx
WRKXWl38/vVJSA9CdDc83/RnoHayQEvstyYVxY0NHVpZLGmRDYgGbPT+W+CHt/8ZG66gbCZSrzJt
AGf5nqLUa5yzVGzWPAhD9jGTsxfdK7abFXCSQoivEhQltbEvs+lfHMDc+Z3lzEJkEjbjk5WxMFud
bjCw62f58pnA8E5ydxQxAlaU2Ve/GeerWsIM2ta1jxGBxJz/APEq1T7TIVbXxyh3iGyvsSdHgVLN
W6m2chtu1ohsRcqdi6RmPIU6z5terVo8Ln2L4RxHmJDwV08fTpennP1jAUAM0idI0KGM3reXk8t+
BxfeoomSQkx1YPXz6N8Hy6H7bhyn4qYFfCZt3psbDb9LtbLQNm8+Srm+GLiQji97PO3OjXw0iJPu
4pJg/AShBq66IO9cHsb87U9T3CEXUh+ybnkElXh9MCPhPSPw6UWoCsAo9DIesBbmbI/AEbfpqqXM
5UxSosteHS//STXIHCBbJ8v/Zt7WwBXtWhEod6EnHbdjUv9DwN4WYF68qWZ1T7IAH7HfXNrJ7S+q
iDa4MkSqIYhon7E7K4wC3cnR2YFQLKaaRAvRNBDhRumELnZg07S0xveOpYxs/3SoF0T7KbhDxVor
Ohh/HfkfcY7WbXmz2RFBe6daGnoCb3H8zx4+4jO8bqkSy3duoNhn14+3AomkKCUkyC2cae5bG+qR
BH1VH6lolpbu4vHhbmser0Nf5uWnVXjKzQQPJUFo3I/Nxt+fUU0sBXfv8kNHzNIIuRuodR8RODDw
XzueLyAwnUVVVO4HOiiayJxh9p4WyEdBS8Ofs0KZ+lavfVCaW81BN6/DV0tpha4bwEbKuWv61Sdt
2Sz/UqeAl7kLj4kE14RfNd1XNHWuAYkGi+7BJppJSdl1plvfho2hOAcQyidh3n9HU/rzRBGRFFKo
cpZ0nVg9k3UlzvBp5jrkheM3duE4Gp2yAwCoZz/3ysg4UysDZKQkUKqJ35GPl/uq5MO+Gl1jUIjK
SEOQU9CctUWRX7zypJmTXL9eA9/ns65XHnIiK3qe3Bij25r4WI8JN1SILqXCB0E/TtG5CaLDwjKn
a1lf8JIjoEPKstWp29cBVBbSiGgokZAdInhA+Yw+MtNmGu/MNuwRGIvOrSmkx0egIehIc7lno4CW
fQuIKHL6G4uL66UlP5/QNCMu/wbGLitajYwxxRKRuZatupmS24h6IQYRVCm7zhwROQ1aoptvBm1P
tlHPoN5TdHMxQ/BYg+20I3wLAmtnDLAcllBMtu8oCwBLABm+bZDBYTsB8PRDbOUZB5aePn7DFftC
N8sspV/6gPYrqgBxhy+m8aWS1Lp/ZlS3nFfM82bzDK78Jq6wjpqehz+qgnrKFmrX1pK0dlt13PdJ
BOifXvK92ggePnQlXqLdNbuICMYWg5NVFaIWSqT/4QoqR3UJnmveFD7t5mJk9B9NreuUt1+PYCQh
YGhuiDZBFZ1yiizi5gCgH+pnxnTAGz2yq2ds0UyFadiCDut5XlTUsH19CelXSQ/swzrrNfL40A2W
lm2QEg8dRLv3mYaIiTAK5z9F2UWfH9NTPmEDG4UNPUnPAAX9uQLmKN/lcTpOHgTU8RAMkmnP+IWE
35RuJf3slD2+zpQguxxMzv+dETHX6E5IB6weC6rI5etqdnfet7ji/B03jam2AJ9aPozBz68F0daP
dktIFI6QrjuR6Ah84CzYeA8CFYeHIVocSoTJhCoFux5uvul7SRt4kCJXojYIF5BcsxvNc/1+SFq3
6Yq4PPyNUnqu2zC2HPQCIlRqQJ9n+DENO+UCX5cc0Kuyuw2WBLVSc5fWHg/S+nQqf/ox79h0yBOD
PgwhUUcy6K+wGs6S4EZsZv4FW2eTGeek1XXPyVWKh+JVUeJrjprIYqWvq9RHNJ3/PvNclg05bVIw
MSjYJYKZkmBC6qluOfoMUmd/3rceB3Kn7ZhzMB6b1c2J+2iKsmW97OENizj/1AF3EUIf5beNBvBL
lcb2ajX+KLZEcAt3OpkpEYpAjZqvzmf4ixTNUXEzA/1lxb0NnQG3xxJhvoanqyvRDXBDn2JngAuJ
24LSHTrKPe3Q3Gro2blMU1K2RhvxdxHxZpAJuv1y3BykaDytji3gRQUdW5icg5siONDvptjijkjn
J+mTbwZclbc9Yxk9+fCebZcpl8+0t8ArMuKinCISDuuz5MUti1GNcfGGqjsCHDYjK/2WbzcQPDWg
IZzdX2vRRgF8YNEHIOB+l3ymtCo9pbLBoMeG1gZOYDslC9/vCzVi6D1DBh3NSXlrBHr2Ey2L1S+H
GNruoImd/NPmo6Wl6D2NIc8BZVH/tzBV4CV35AMgJ9zr4QiluhHNGpi4ICJ2hLJsR+tQQ0NKLs16
wn4srA38N6D7lqIL46Y9R+vQ2mUQXjvrU8KhMBcfzphNrn3Ho+XBqeMzvjoAB49Vu/AUqhboxvqI
Zp3oVRCm4ywYbCmW/hqjw3GP5vskzobF55fVTAHRC0LmMTOWbeXMHQhqDyrr+GVfkFmZaN/hx7//
Qe1dP4JMlqBwDkeBV9WSIJTYfI1BjSxBqnXF92EAy21Os4gQdKv6NE1WKP0TLW5EsEhToRDmt4Cn
xT3iignXxgeozHo5ta/zS4+RIeD4gr8Z877Jkb9AY3xpdoPDxJdv6YlhzOVpmaTf40N0Akxg8jjo
ts71O9BWUZrXqVShYKbdFqx3fE4daJDkskZZC4Sy48eGQWd1aRJIx3qUm9oE1VNPPlIJjRXh3Wkv
flREWefiZC2r3Kg7Yn8Mo+T3LWVkAcPs5QFxC4Dipq29vayv/WtdwTvH0fAKqLikq90z9IPRr6GF
yvtOIGGBEQQQEr/MJsBdNhINSguZ01dGF/OXeIXclkHnlO5lPI5pGGCCEFjuzoCbD7ahxJ+dTTjz
xoKHEmEeeIrcHPVCe5TrG1R58eG2ktiCaMg7nXnDtezYHzH3vJt/rvHwmRFU4G6dWtr9eSY6qae+
Rt8vO2NE8IkE3CR6T7cyYK8Vtntf3Xm05YJX6nZbd+DBqa/rYFAmi3UulGRyBjZbz2Bn40T5BQ92
mEyXBYJbEzDZZsDPDmGMC4QkRTo4DxTVlkF/zb2usp3oeqbc/iQxHaSgiHfHdowgwUngI5snJpp5
pacrjnNq0wiEcJgwxzGbfzZWOZFCoI1WA6HIj++BH5ZFF7mu3zQdai+ZnHkgiFtz8xD/9Z1ENY78
nJYWmb2F22ez56BnSw8v6s8XPeiwCUFPr3jppE3Ncx+2WXKtK2xjaOZlSWpJRYt1Wa/jBuewH7tQ
f1JQA+P0siWAYHFqxAdOt6sHl9F2YSMen+eFjxJ2nkLwCdgePN5TkCVF0OjprHKk4WwDYG6v+8El
Y5uHldXgp0Px5+uv/TyuxEp9M+w0Vkl9hYY/3VFAq0EAKg9M/L5gN+5u2cvlF8kTXPqEKiiltE1l
GnhkZPL9ZUuE+YSrYD4c5u1+50b+o14XU0EkYojXIwDS15BG1wugvzH/R7CBuzxNtrzflVJ5NB+P
JN44nxMxlg3qmVlKAcRV21Tw/1SP1fxs4XQsJlhw0yV8+hAIQb99D7PUZXnW/PuGqKA5o+KggOX0
4+O6kYKh3JIjWn158Z4VafcuKyEdRYjZ7IwaoizXcBHSarCnJ+IzAW8kx7MXGSiW6X1BI47hisnj
bbsgh8haWlqOPLLrTcejsunwy3EGnmrB4c3ULP0mmBUkxIN/DUwgzQOWKmepvEBVNaBgEB66XaUW
Bp9Z/3Gac+9jy1SZAsF3mAbNfSJQE9Ti1srV7rQuIKqfgoEXbXzBJNNB/q97JZ4AzaG3vXyl3ofq
aKiaIoI+ZfSKAENY7N/FdiNwmUuyMSbC4KZ6l8evR4DNxP6QEWZKnXqeemsyQdGKntOSEK4f1j8f
q/PAYAHd/cc/swcdJ+jpnC3sSNScjQCPtY/uIkULC6bxN6hr9OlviCjyWc7TdUyR7o8P/B0ZXJfj
pYap4+ahFS2UGKuo3YchdrZwlSalvGnh/x4beFuZJzrGREDh+/jAtt/norW6h0xw0FosMOwwh5hX
gEp7VPk4VmBfAu4sBh8mWHjMF+4mmPvZJ1HReZeKHqB5ETCuhTo107UE/5dQjVY9Rma1Y2gptKF+
+MSjM9ApVjmoJS9goiIuoBWYwu0u+Xo07eZcE0xc9u83X+w4PEiqRZXHkwtiteTTnXztQHHMoalK
HgcA+RsN0i3TJapP8iWOfLKkRgfKNfGJYiCoRpLdq06DkmE8o7mWUui7D+ViBJ9v6G4ovu3byoeX
cBdhGg0wSRvUnrVinleYmuSsou+FUJ72tZG5EvMA0fci2wNESEosP9Ld9tlF/WWaM5Gb7psqbIKq
IeKwIFbsGkusIxx+sSFkekw586mHLDGeH0icDt/GGHOvoWe4pAb50H91zZKanLC3h0399cx8PDiv
ameQZHLUPlzuv1FEmeMRN7a5SnsTL9JPMXVZBjBizzJ1IhU0XTs3ADVYPp0ufrLJ+sauCkJhx8tY
aZ7sw2EkMB+jztlvhyUXEtFcG6K6kdU6r1aziLf4fIFkoMQGDIVGRAikjylhs4v4Qixr0S5J3v7X
YH029YrBQ4cDx5mZE5u8Z/9DRUdO8sVDNGxc3nYXq+wlPGtk6a27ecYgLOcCPluM66aC1W/dSAUy
gG424UxpDL/MA1QxQZADUxB311FwKn7yYd9PfuvhBPF9D0S278KqY58dL7qGJqwnvRybZXA09sNS
lokliY8WOMwc6DcsqE3fFCitCw+ctOVGTFjXfFHkpy4yGXCXLImZS9OegWMrVic5OnROmhf4Cw5s
/lOmTzjAh+9WvASdNjT4y8d+4cFlCGQmOo3STjm3Uz321Mp5gbrHSnxDgohV2Ze2HsSmMXcdFsGx
uDkKSlTbb289IrlMcQy3kj7WG9zBwZCSf9GKkj8zSjwET0vSNzyt0cr5qdQ6ZEILT4dDMD8lK2oU
pDx/96+DU47qH6jewI8i/Hr4vH4bslmU/5P16CyJbjG2g49QwJyh8JwjMuPyB7cLA+Zq+LRajkPV
fasWD4ji0woDIj5YY9juwqBoVh+SfAM/1sJcVXd8+tVVykBG4p0OUsqsuRzGygE6+W5uH47Oqc9e
9QjuGqHBBYROeNXy2RoJsnl/BOtRgBOCHR7RDXEsoeWXN5ozLBmUAFGqa0DQXzs1kGaKdJAl8A06
cAttLoWvg8qw+EpnSXf9yg+FuyNtvNEDZm5OMej3ryq5asuvmeNsIT4mOSeUztYclpLR1cZpuAZO
uC75SD6ozDJdU9Bfh+5Jc8uP62TKnTQPqc2hksPSNI1FcgTW8sXrNgVpiDKECtwmLFx2YBITDSCd
0A6BU+xls+lvV28EG6jrQDxbURfAMjYVJCOSdz9hgKlvUNrC+MB9yXD9qLUF9JA5Mmyvb2TIHAkS
RwPFtARrHBSBEybo2tn7tG855LOI5Tycco2tM5zybLS5fv7J00AfZYW2tUtvFsOr1N7lifutkFCd
XhXsjlljv9nlsrDbgASqw/sq4gFeQfGmCVs9K5Ddv/Yq6zIdTrO865E7gKNiS17ucVOTpMRNXz7f
C99Z+07vCIVyCNHmzZpW7PyXx+joGaHta9eDyjudk9dbym8u7R5ZLw2WA4e+RplXXbnh5u1BPJ3o
pnZbWD+uk+cnqaLl2740SI1fjxUuh2kS8iL/UuoolBL794P0CZ2hvzrAdqb+Lwra5NsvdHfc1ZtX
ySUWEWQl/vOTPhaE2jaoAZll+iA9NdGs2SHxEN06m2hFfa1fElc5PU0XvlAu2pIdhiVOzzpUFCNh
/JA6AIc7fgS8Qp+ZbRowKiUCgX6EuO/kcLyx0GXgsa0UenzVmHBIP27O7nEQuAB8zNElACErw4WF
yT7/eWDduxuk1mFQuZMomggd+6ijmFZDCP1poTO5wrmXSx6jYm2+guwvKkVbxm+tEr/5l1KON9am
CgbLPY86jVo168soIoKJGo4N4/W+Jo1weY3On9e6Vgy5vOjPXFlndlf0h0dTZLn2Ae2xnTNM3ySG
PFyBbgz26SbpXkkk+wW06YTIpB91GhkdzcK0TQxcCdVWlPJI94ex/ag8a1CvdMXLDb4WW8OcpbFf
4Gds1nFHetCAfVGGCivvutKxdfH/yadhIXagpXHEp86gPCPklMV0jQxtfTf9KidHm4QT3nyzjJlQ
0r7HYhuUyiy9I/7++K+PfJknHmqD5r4cMZ3S04TKtbdUZFLW+0U01sfZ0+2wTZDVq/jpysYwqKuZ
AOTBQ+2mPDJ6WHVw3gUh8RC1X3BaYGQGZE0gbwWIKg/QXgmqcmVALRwaag3+1Qs7ZVoxlWx8zGD6
r9ew/AQydoSw6mzErFbzrpHGB98ZvBHuIw3kw7gS9Q87Cxvah93y8C5uCw3qxfKuIKKb+W94kORL
vyeepxm/8BX95543LJM3+qkvIOZLlda4cZSJd2vO6pPTzT1yH6p9gZXQ+Zn886vMuowTBdiaWVqy
Pt9QR1Oih0UwmOP6AIa0k2auLOiKRTl9HwvSRf0ryyy+3B0WLts8six6QPI82V1OTEAh8hbZODJ+
1FkDJonyh/pehw6DgAMYZttPOUEZMOYSix0IzdDU6reT9DgmI5eq6hQqR0KQvqWbR2WEck5IZANQ
zt0hhdvkXAZyqGOWbCpTfqG3kVG0KcpViUsZ3vtmE5ElT3+ozoNxSgZKjufy+vYZauGjOyrMGvkP
lFjEkmjaMp1Os3buQ0TfvVaDDP40r61g8d04EKnBYShujj4zjD3odhVy+H9dQ74aQDCHsNPcxE8o
/JDxKh/OexlkKLsfQ8AhLMKEj2Ir4i/ck1VlN4hau+WAX39i+cYzRVhv0GYoIhJ/R9yauDxUbf7O
BewbzmP52HgTGx694HsIGAx2y08vq2Be47fGxN6sOi6dmZ9ndZp7wj4Mh5K+Bu4ZDbSjmBZ/qOpV
IllOvxaqLBQmZgH/H/LJAlT02SVWAfePNjE6soyR+iiZxezTOcGNccF5nmGmdGbHVhtF0LXB5Rix
XJBU0Qbaqtnca2XKVFoTIs/UUXKEUpjeKfQQxGtbKhIto48i9nlCZWWUEqQjFsdQXsZJB2qAWY9/
uMRK3054Li+tQJwSyMYnDFETdpjZAmClHbd2sGyLr20rEAhWqfjJSR2u3DTkUtC3nhPwrNF44pzn
S2Z/lyIZvDb3btvpuXKh88EzXWisvH+tG2/hwC2WijHeV5vpuF1yggTaxNmrKOBrZq0ni743LP0s
v0bscsT9ETxxvWZnUGVwuDm8MLcUiRss8NnmEQ9M7+sbNZCgzZ0+CyhwWG5G+vCLnGFKwb6Oyi4H
e1nlZiouSgzveJ6RKXKEgtlPL1CJSKXsPHu7vd2AEZ9WycVY4urQniq+yy9JCp1oGaZErqQ+tlQT
4yiChcuuSCOFlya4Fy/rlkdaBZPYx9KOATxX5UYcTw+1RADNePIUXCweTvGMbnNdlb8apdyddmO2
sMQu1UPbasjW2aoZw6GOWnrBfryK8Ue8++ZWV1aapFf4BMm7UuG8Vn9AbYKb6U4VBvUE7uxeuRq4
6SsjxKmqBEo9Lpvt3xBm6FjesOWZwz40kn0tfBgjQEfByA2aZwvAxA4jAiYwiSQ+DjWX0N8tdyBe
8XXFu3lcz2aPBJxT3U1StSD+TcTiXohc1yoVKx75gVeguSEt0hUZMOWWH1qz22KHvOOdnSumwnyf
3Fs05Z16VE6vY9zw514CFbW09KD07cA9TQSxul4QMXgWxhpdm5FW7QgSi8MjWYKvMFJ2mQHz6l8Z
e0B435RazzA7hsvVYsFJ3cUUa8ZiR7VIMz0O8/ZWsPuqia9BDa2RX7xSsghLlVN/xAg8QKcglffO
iJWlTbRsNBhuh+utscNE6SjQDh8dH6ZiUy8S+s0FqTIL4NdiqCj0q6JIlcgW9qdA9BUfJ8QETLSd
0Pkrd238ekk2P9cCZqG6l5iWFgP/DsYCwbtugbqlebPphh+qslNAmLqsKJ6w25PCEGVCQA580XyA
EA8Lju2ueNW2prah3dNR5retlO6oOzzV2eqIhjURQL5tylgunABAfIWdJ2cH6H/8+rXNhIeipaCn
ST2Yr6EcY5/Ny6dHsQdnCr2LGCzwmEFbtpkZEmcfYfVNIZAHkg5MrM6WKBBj1i6DVM3oIVHISD84
jIHZBydy9yMD+tTl4LcMNyEAsBsBM2kG/RbhuXZdgb8rtqQaAfFhLgKCPvVBfTmGNz//9PsDnsg8
roOIK8xmsnY7c0HVZZ33hZtp9Go9hj4YxscspxvcL5z1UFBcwIbqNsMNUYonnPdiGq6ObBVwITm8
Ou+5eXf00LA1lRtsqycNFKzef90jue7xdL+rTpFSt5Mc5khi9b0fSmwJ017hfZcFezll+5pjpy6n
liFpyRT+r1brO6ns2H4LEJMupfxV8fGo9zSDKeuWGP21zb+x+1CywimE1reTM6H27PsxSQ8NXf9r
EtOn1A6rZJWmmKkBz/cuKa7yZrkidfuOMHYA3/Tfjhga6aAssj+pPAVoPlEMJJryp0z+5NO/pDC2
HG7czwlI1B/6+DkRSi7pZQmOburh2zZK80jm+E0Yccouad6u+dV4Is6Qm46GdGB98HTNceo1/txd
1eyS5IimaFDb9XV2vQlYLKXnDjH+Bxh4rzNGEiYhwB0u6sLhQWZK6Y6134z0vYf0d8oNlXK8YfbT
HIFrR9AsIIGyntEXelzijnHC1yr7Wm0EgMXW7Pnt5mW4dg5yFOR/tDfYvOr3cFUOdRd8qkIZtlRd
p44VJXR6QETzsMBM6D2pcHPK4lD9NuYfhjAJoakw3XdLgipSTCeBlh+uwv0hReV9G8o+VeKzaSZx
/m9ZKnbvnmK20U/B2U4wHdQj/E+JrR+K43FtUu1PFvdxhRP2NgCZoeY7ZjGftnIMMwlgVuwciXvy
Bf0fZNSyms577ZzjtUv4x1oGHAz39hpFJlSf4BeVibms8otOpobfnEJgNIK/WJZKUeNILB5+DG4L
h/mAwPz2re42pak7X/NlDQI6efgrM/3Y4CYeyJWM2ldX3NX9Tee6t38jH856bQbdx0dtSJNy2uop
ViiSb8ahM9u24PM1OeHLiGjxAvZus8oS0qZPgsq1UF4z2jJd8VCeQDVKWOHEO0Iss4NWQ+AFPMQV
EYTd0Qa/vUPY51ma43WLIndJCfgsI9FZMqpcULD5DeZkiq862FDEJ8Jcu+AvBkGbJuj7MObiYIGo
t8mqay1vhFx9tcNbZSp0rGu3x02SwxZTNlxjD041G6TVWV/S51qWhhdPiHSGIRvgYaeRazfbWse2
IFi3Se7GToP8jSDzBBHN8Os8v/0pCMgYKn4HGSJbcRRM3FQySjDFPwxB/2E5PqBskEn8mLYHDS0J
47KFXBLmGF24t6jtfz/98Lb1t4QPSxZrr8MyIgAUoK+qkEiS+vut+ExMJy6vpmVT538K49arTVks
modHb/6MK+jWmDNA01AtkNbnjnrJj5hcbJN3FydZK8O9HJ32iKhrgoOVAWX048kxxgfc7NwvvtYE
zyBAawphQDOerFQwtGBCL81L7oAmgovrGRmWGJZ8fbhVRz3OmyNpEMijBiA4b7+K82KqI0IyEgw9
Md28yxIzIec6jKQjeYTfZKuaY8zI609Sr2Nx65wV3l9u0qX71k92YMMAf012hq3YtRRzoERMvxpg
uuBhPje7tx9Uu/9oIF+NXO7ndrXfAfHgiC7C97hTRRZNQgw3Dt2uScSmhEhTetz3OU5vrrIpKcI+
QXP6MU+ozcWlJbaStbqTQxS2NrjHh+C4R9nOAFa9WcxNqnRt19YjnGlnSEw60K/3266FEEeFvHoS
kW7fh2hSOYD0U/pIQVzmiJtTuxGrx/K8KCZR8EfneVsiTp3DKGP3XDVW/9ipqfRelAFdvKaCzoBo
JhyhbUaEYwHP/YroJwg86Ac43i+ssAeWO5k3zlMn+85QBWjr00u61BaSHJk8a42kr50AfhqhzuDJ
oS/MKwweCUbILR7dvK/6LycfdmXj93JdrqwT+h0Pw24r8YHkYmY/5yRSziPg6jNYM7f8fqFEX4v5
dSoCx34YyI2lo/QIBHu6he0J+Fg+LWGxpv9eDyYWK46qCiUegk0gJ2ispm+946qW+liEGDBVTtQB
lqxaD9ZDZy55B9ZLiB1zO55KT+ls1WRYdS8YD6bRbNRN+Mlc8DlIgEheuWjM+GpBtvdCP2I8Ieo/
tBz/sWfFYIfrtj1pJO2zL9W11gw6oOY4tAwbdjrwyBE8UJd7AJGrhbOAQpZPUQVrxeWP92sNJyer
BkoryKpVQRv1LOmIxFi6AhgaRDngqhYhA5nAglxJsS46Rlr27TqWlsU/gofKfnpb3sLejxZAlcL7
cfEnckF0srj6CTARKVS5zLIbKk1ocUnmAxoJkr98VLQ+buOTwck/AczBW/JPCDhq7ibaW9iy0fF9
jHfX7s5+vOAct9dBCYMTdegdpQctVxOpuKHj+hHBmWx1Tf4faE5ccTC7dKAtmk/A9j3kVhPRZxnI
XROlPwRYvXq1o4TG3ggzCxKHcp0r25ze+8siOkUtHoL0dewr1XOuQqgPsjUb3172x/zgPNGKxAka
eD7alJ++SA1LkpvJgzY/YRGgmzgkWVOeeHcNtITSsgirpTaJAJ6le1bcPIyrg9+BU9ZOQU/OpyXP
JuxbhCJ2nyGxsGbhNry6tobV72+lhjt2lsxn8FUdYP0imFT89QXtuiyu4/I3J1RvtPtu8hFaKc61
XDq6OmFRGw27mHaD1WDAwTlbib1/81cbpm/DfnIweHgkXeamuEoQesQ3vgyylaf6VXNThovKcfbp
hmidu5elSMJOGwf6rVPubrcLqRojyJTP0zpeb9tFr2el2NH41jJHgnmBYsjj5MBUjctexdwbgymu
PZQ9p8HuFpvC11sB0GkIbOgF+ol4Ecg0PGb8fZvQqIR1NFZ9bLXe42Em343vGks+viU0NvNA9/R3
Un1ycaCgQKOrR2qcegij9Cf0TIdppyE5pQGXYxy1J/9PeSTA0LHlhViLzg3myasXJm8S4xO/3urg
QZmfFRHa3HoTwKDXNHlQyq2GlEBHDdDBeKsETPgGwo7bKKPU4fP+L/p9KCy1LOQ1by/iOSmYvG8u
ax89/WtTVtbCRupWo9/U0RXOwMNgU7DHx+4RuEWP6DC8ODChk5nNq9LpjwBp67Qx3k1l+KGMsSBc
MdbPBQwdH4ZFMRcyDfhnT9noXGHqrABprv9S2qKeTucYzYD1t34ZK6DCgFFWR/tZ6oc4xS+sPQ6i
j48LKsUNQ5qmnq+8HY24sg28QvDqbp6B5g28TxQwt7g5nPW17f/OQkzkEm6zL7yWYL90RTvOroiM
zyTE7ad9IQz+JM7dhRhmen0YNg1vCunjRhd4S119mzFkRQ9iCQei6MDO0DbP/g3nMp2O8bNVaWmB
NfGf2ZbLsXfGO5cqLho+aqP/B4SovblJQCBiPpDBicUAqiAb6R6LBnSREH76qVDn3aYXj5hMYO8J
ug7Zhhrwdfl3hDVH8Gwt6TomZOji6TcvYd8J6JFqhwhKK17ruJc0sPTgZsC7vevCZXSZAv8922/Z
Ea/PO8+2NuhCIKnZgvYoCkUP1PuuGH/rg69BToQkZNV2X3RMAvg99e6Ioxr0HjUnNs0MJe/t+8JX
cIHCI7Jutitjmc9XjLzXhhBnV3IH/Mh3T+Srfxgn/zI4pQVtitlxe8FBSx/E4xtPowHRRNmJqeaM
6PIODROuI4hmIVToNVYDUnVDFQq/cRft1IYMSZKX0yNqm81LIQxiHKHUegxs6PjBHN7VKyer65nz
wEQcFFG2Ra45W256KL8Gw2v+33fEjtq+2rgAXU0enazW2auWD35U4jSGqMRf2SxPxsxiKRbw30Jw
7W1AQVJiOz7oq/L1uuzL3nrgp50YOkHTpf3IQEG8rvIdQRgInSXe1En3azLnas6MWpCeybs4bIX4
m/XKSQXQQC1Evrb25QOfuzO3eGxwPlLpLOcKrHTeeBQ+FB5qKtnB38gBzpovz18Gz0gUCPYqIBpK
wF67F+yrUqeCfJQfvBGYJE9m0ikKvOTNHM5prwyc58ixGYqvBbsa4V6ajtsM0qQXcnJX+nSeRQ7Y
clS1qu+qqWylAvNA6atFGZCPhDFHDCLTEhW8n07SYYPHf6hkZjkjMSIzVORhbcQem8Y/4K+QOfCk
EUKrjGiSz9wdFLDaIw/pR2SqV+kmJfhysg/5Z/DV2HMp6n5EUEkhAkEOnUPkdo7nXlUgDdbSwvtc
YqaK9UtRo22FhYj1zDKDLv1u4noqVoiJXP5MealmEJkWJTUHjny3yVzPK511ceTExG6jgyrX90Nf
LSCwj2rFm17QTxjXXVr0N3ZhcL9nkrSJCkxLF1294QFB33mRH+oUckL9lzVVY41s5uyRCurzv5/m
QQ+JpyBy6zWQ+NSqCbC0yBtnv41W9jy61OecXXvs3d7D0ReHEo5QqgI0iZrmkRoVvLHKxjO32eCq
QFCgxbObpCz1na2c9GKt40hboK7Ikt9Pxkej7q3kbg6piSp7hCmsaXTS1vru9pAXelATK72tuCcJ
eiymO+WZgcNAn45xPsdR3skkshswqGLXvvVyqSf1SmYqdSza+M/Jlxq310gMtmNO/iTJ+HTl9vE4
9Tc4MZ0O2b10mguaDIBr7g1LyvuWUZomOiHzIwCmCtsKaOT2nyX5Jn6mchN2LHnMKAXSiDgc8hTa
qsBTQgLodTD3033b071u8iTBTpIiESNpqPx/LqylwPh6uT9FJsYZ3rubbV51GXMU2RTDsCVYlSyw
FEGDAsvpf6L2iIqyARLVYCp/Q7KUL/A4cm0gG2Fzf6UtICfUGjwp5dPoKqZ14pMso532jXQnC0N5
3u+XP1yxLcoW/jVkKTIscAlI+THhHOSQBVPSGLqusP1n2zqEFMh8JZE65OuzpN/NSyNv03epryxq
gIGxhFpG9MkRxUQEiUPM1rrTCGW+rNBcVHqdrXPIrSGOBEocK3m/jxyN2EKadu4AOn7IDP145lqe
VNpgzkT7alvnzFPssRyg9kmIhKzV0UtbZDEFmaX/hHO9bnUkWm4FP6RU4skaPB3zTTBIjM6eKzFX
h8AHpSUSMWBAIT3jHYGTTqdwf9NeEgTL2+uFmANwftTH8E/1Y9FQlmGeMx1xT/1Vd4p0gAC6Bx2L
xmiapS92INtk3IfKu3S2e8ZW7f+boMLwm0QT2SEmK3kyn9Wg2vGTyPgseI77G/azVInE073z91kh
gKnLj5JD3dAIL1NJksvGUA936hNBnK5tX6VY93sLa+33FSCqrWfRl/gLp2+sp5cqiAbn0LtlhJSo
1NkMW7sTOU0E00yc5wlBI0Iwh+wzzcoRQzGlGDx4/hjS0HFNPremkXLA44v+SOL10MyIggnbPDZ9
MRqrXRFgEVXAbhSFzRmti9hXa6lqEg2uXKvAriUaVG74CRJxhwoXK9KiZIDigGO5+z0jC/DtrQrk
MNheXt+UiG/Ry5WGUl/Re/LnwEzM7i9Jgfv+evSxSyktqdEdEC/HhiM1cEpmTxP0JEkgmb74aRQ8
iQOWAYA0aJZebGYrSWjwL0RUOtQUfR66rQ/ZuvGaBfFL0iT/mEM8J+6oEgbgtID/MEFcWMaizlUB
ar/t/ld/nO6Fxiap6BBiwH61Z0mieuvXrXQcac5QJTjFMCh84IQPauhztF5FpPVweEcGGio5wsTF
nryRuQ6mD/GIQnVrl1ypZ2FV5RDmOA7MAttmpvhtO9cX7aLmBg04i2xva0itgcRsyyR3POvwFYYq
A1hFsOD0Y9Hib75cVsaHmLEMaUJqkLyOVI+VIktTwIDj9Ec9aRzdSnbIAa4cAIQ7iDrQPhJIlTO1
hwOW6IhDjqOaQVBkTRI1oTaL2g8ZiEagSTRwtWCnyr+Hcxeg11ZnmxO53RyoN+IYuzE8izysfgbS
1gEEd1dOL7VLuwdeXFVvUC/waybrWogAJvQDzrgr2iiW1EEOj3hwvItpYExcbwa5jLw4hkAgFL05
3oqlnXiDcnqQj6mdqXQK5BgLcYTziNP7U0lCeH9QseBFsivys4m0Xlha2PmpcGJvg+kRu5Qlvlrv
SICAu9476fjqR85NHRTGv13rlYgANSiQ4xlTDVNze2b0D3AY4MpH/rQykWX3NkNcGhahBKc1QIfx
3SoLi6aOGA4CeRUXs+SQ7u4MozvDkckBnhGBGZ2Y78x5gfVG9D20DsBTgXxI/iRSUR1O/paF8oiK
yF14XOO87mzQ6DWKPoxI27L7xIY2v7Tx9ySUJURfo3b8MCmeWncxjB/TKBlpURW6SYdWskEtWDZw
sKnZr28DqZRWHOTvJvSbkXYhcVGWSBod8vCRdcVz+6RaLkl4vPYHgEI2R2x8pMHVY/BaNoEt0CWh
5/gJSLbh+u2AFrqkEv6ZI4LjOa2BOtmsbIrEA+nYWfPczunVoSPo7XDUrD3J6uPsrbfOCydfa5bp
SPEtk4dZ9Ene5uNZjyJ3W8PRgKvw401aKLB5s09IeLnobVpkRbBBYHUy3V7Lq8SRB3AYT80q1feZ
RTWN2gakI56dbukVTtIH30pcOd5WBmVO1NVJNSf77AXbT/2Uahey1TRrnr6PQyDpzMlR5wWunBQi
W7zVR1oGfFrIF/+9C0JBgHfFyfb1N8lWN1DQLwZda55kfY2LdMitr6KFpauqqM/hc7x/+FcZkmA3
RoGSS4rSEuF1qkQxOsF3FAujS0fGmI3kI7AWpk721+ZlnlszXlCyCDEVP++/TKtfeYhCHEAU6R+W
oNb0YIU65kZdTtiMDaAXwhhQ1UA/S7rDSvVgBa8kFTEyCgKdT4sXPwdadz4t7ioUYPjLN/k3VpR+
h10QYy2dIpzXhj/K5pTwP8kazOjU8RSKcpBGDdgm4GfuBadcOXBoLXh4JUBFMU7HstsqPagRhOKZ
bKc0YsZ/JNtGgGiFTqUvN149GheQVFV42G26nHD+gUSHw2ckM5s6sbDsCqHBW769T1k41zMmSHLm
WpzLBPEoWq0PaVan2P1E9CYM/dqXsFL4wbZLxeXOrYfgYiGriLmH0gPqAy2LwTIZo08kU8n9bd2H
9Z4Zfi01XaM1rH8+uYSGd4oj6DkUGSPkLA6ggHySOskcekGrl7LU4LdU/RGSw+4J/x2+pPS/Y1dm
BLgjUqHz3QsMKaVNtYCjVG7vJ6UlEnlZsLIN/rSMmOaTWjidhI+Bl8y1HHUv/ntlt9wjE/4+Z4Pw
afWhu6BBwQm3nqfl42TQbwhrhtDLIjOJBkTMIYjdwOVPnkdqMZQ4tsSzilS2uPFMXiggnIei6KEd
oS4O/SO1PjhawHoZWxIS7h7u9wt7tMAcRDAfEmmvzphaLRIBpJDDmra6ODopbcpL7luWGdJtGy0Y
gWz2+DzPEnzMqdUjLd11yJOJ5d2NQZfekq6GSYkFcQURD2eJw5lf/CpKpNVFwTU2EdrbbWNuvtWc
xw8XG9oQI6tDE1xbW/05p9oAwJeMvaTlyhOaafF8SUzDZWgZJ5XjWpQxCHmjurHbJG+ShuWCv2jS
i0Um+/GYIYzphq0CFk8A3HlfVSPdGWYHr24USIvsm9z3AncsRsduW8di5dn2UG76e7duRPnIuwqO
r9fZQax89NhuB9HIa2UF2O8lfgjtZIaDTiQOaNnV35qgzs1oDMKaIq/WeA3NWKb3UrcaG5JNCiF1
hA30hCNLtkogrr4KxYjNH6OSkjrrdYawedr6tsTvOhnabniFomUoDWgD8+JqnONVYg2ocHwx//Ac
kqvYjdMNrCkZUN6aPmxeqX69WsqhMs5uML7VDxYPeJOuDAXr/wieotBEmkLCl7lMyCWSB95+QKn0
EpQ7bj+FGhJwzSu4DdeiPP3xWqA+4btRfvbuFpDK4NXH4YEWNVdDanaqCaT5Esx30smKoSHh4ZRV
2xxLYrMaGooQtcgR7v03Le9juIry+XmB9iirtb5Ok1JrW3OvYZdca/6CBli6csLRkXV9/U5wC9w+
8XaGFOU87fEBhd7ACp6rLpwEVW+AJsATfBWf2fWFnz+oBPgD9fLqBFDYP+ijfnhWhK/jqlfxmA7J
TnJK9FScQ4q7QBcM+EcMnR/LAJbrtIiQcoLRnxnGjdBYHpmsSWcKIXdkWrmyVYrH2lULLeOmFB+R
ReJjxNX0g1Q9nKarpZze3n0FaNASsiVByDvkPRjMSvYt8lAXHES2c7aUHL/9+qsej9bMiraHvlM/
0Nvbfooo+tl6+s0vx8qVhQ3X9FhFe+hYXMwXq9MUtm9umRGQYVEQnbUscf3pvvfZXW7t8zDkJoWu
vs4UPxjQB2swvdrnBHCOaD+RYHlEhDj7ivhb+djkl8GfVaw+jRz7PIwvNkLiJThHFGCjEhp4+ScY
7ciikO5hX/xgi5TFp1/iJYF9IyKW2drwEprO2JWEv4OEBRYdhRI3OxZ33PfOSgcVewHaFzLYYFlY
3p6GfjTvKcJsdaAaIoMOuuwlnEAGf3qoCxADpVFBCp9UgWe/OZWSy+cmxDokJ0KDFhEELvBXOcCU
HbDJAduAzXWrqz4s0QBl8PLrp3wAfyhZJuWmOdxbNh6AY+xdMaPqNeiiKKiU8GmwBTxdCbmqM8FR
4oAhTBklbiKSdol44pGXRur+JYC9sY3mWR6wHZbVcqUheo0ZCYG+VQ39HIh1r8NB274wdk3tfhhP
d7HMw95JS6pXOicEikLJt5KmCwloriIVevSV25fg/Y7PIs3FUCrSH2BZx8h1haYNBYa6m60UIuGI
Jof2TgbJ4EN+QDx6TI8srFSoHFZPYAhNajrvruDsfw341n9dAqm5GyK4r2q+l5t657Q1KHKcPEXI
pqlHM9IaiFWK4W0kC/2DVLMb0sD/XmQkcZFlxVlEkhI0R+J3AXQfTb2GqFrouzSCKZ0UvjhrERdj
otZod6CnU3mvWyPLldrcs8gMaEqeeerEj5MT/Y3WwoxHmBzUBhrrXEJ20lNoRrJ9QgeuOJOWuy64
48BrrwnnALEvt2EVRPjogi//54ZdhZoY+oto4kgp+JVwLwRZpNRxPDY2/qwi7RfFxo1xceqpxpEk
xaKO7x40CM+QCqeBmTt0nHGfe4PS5JCUZB6hn6y6dpdjs1eBM03mwR+CXGFcqMx0HaPTtQHjmYeQ
RCpCBO5dfRlnq+zCPZdNUijC0nDT1CF4nUxcQSPMLlU47WmKJGTMyZplSnOob8Ssd+Xj6NmCEgl7
eREKuCXAhfA8mQPxmgoQAS6+UpTiVtCtD/wcsdxAFw+VMCYkXpIckFwpdcX0sZ4JLC+pb6Ln7uxY
+/DBS64D/KPMe6KbkL95SjtV6uicYaPt04lM6D35Jrd4Ud4iSeIiM9AIJ9x9Sf+CbaNqdyC6+6py
gO1Wv1tkDf0elvF7HQVCC1/8qyYsIOyuQVeE1+7g9YJDMhjxI7DfSVIeulKQD2u5OyKpOD3ou/Q2
jOo3LzsI6Gxy4L4hQLb5hHFwiveTWjN8CfvaawbhzDTUcEGm2bpH3dCjGzP7jeROjmGAE4qo06+4
neJpti/TyuCOdf8R9tDkHID5yNW4e+ig8EapeKVR1M42YpMglupyQFShGEyxZPlT6rz6s4Q4bcj5
C5T36Ob4mZqD6yTThtuEX+E9nuJjPia6faWbWlaWbNffBnZcE2ldO2KVG4XPPHgGhhpeV/V0Njzr
lQri8B/EyvckcvRlgl3A0tETcKfTcOA0j7AsRm9M6QfXfRV6PkfZSOEkRlTbtwgVFrucz7ZJCUh2
iEZmawiLNfoHJI2D4kcfDDuEE1EkEsokPEiNRhJxOhFurLEQeu8ISrBoCOrzkcWTO3rNNstJmZoV
m5adNg9WAWIMEfEjGXiuTLmd43rrLHtFBbzYoe0ubzbecpgU5mMGiD6pakMQ+FtAd1X+JjQpXQ3l
ztY5/MYkfk3lxlLKsbbsBHyPXVed+3dbFJ+zEISHu+9amKwCIQ9J/E35QWcMdeRgv45nM8qHPpdk
UHtOFCb1B/DZm5OgLNtdl3lM5osGUsnsiI5PSIRGRxgR/W7GjmkYJGE/4QI3NLmuMhkBPv7jI/vc
uJ4fk9hSFSJHkuMfYIa3afFS7UIFsSme2uaSvr7NiLbQSqr7A6BF8LUECnR//DCApMq9lkE+oThn
cb6G00rKJSy/OCb1d8VIecJCHEEB4b+/+Nwa7o1W0QVX/kMidoUlh/zrEWiS2hvUnAWcv0mEHttL
xwRHbT1xI6ZX0aY9YFkY61V9hIpCJ+x0PR+ZdTJ79e1VmMFjVcK9gOEEJK0E9dPv/OVkHLojeC57
RkUMOY+z8gruv8e6UfczeU143kkpo9ez1T4NdGssEWtHOizqmvOcGyR6EfexUTlEEeyb/GoYCh9e
BmqkBgDirxWbfyOMUiVoE/So7AZ9trIbt0MAoDYZ1wV3y/JU+etaz0Wsz2YtxRzhb9uwDS51DNnf
3mjIdMMx6L2OVy1IYRtEqx5iUBrO/0xmTcZNGpeARBFcAJBuJJb4t/FQu5HmPShX2Az6RqaMJKvq
N77HxfrGEYNNrKKL3w/akg/JY8U5bSogGwzBjimnoReDMqQEDZlrTRqH45Kfr7a8S6NKaeLgDkzd
dd3cS2q21Xh2fJPIbUGX0Ue5ljMwsDhRG2vlyz8XDmDodNbkBuFuzMfcwgOjKRz27G3Ms1h1RXxk
WuXCx3vZj2o2u20wUUR60fpO7I98CAZFFrWOTfBCkYSf85jYFNFGErQyV7LvDkPVDgoMWwzqBNL1
tIxh9Fq+YLozRBiLU5r1XnRMyVVJ+gOrGo/0KBn6g4JOm7QL/C1c14xCDDeUuXcFdbTuWOel/z71
RyK6uZEXtdEgz5/nQm6HLZ6wgy95rGfDJF/y0FddCixM2LHZmtKGDxrGEZpStDF9naTZwo4rA5tn
7QeX5sz5udQcQ+P3QCdYE+FjXDJH+RxBaTmYfaT8hNXFDnhQwxBQs6CNXtmC7IGhs3kPw8p9Fagm
VPWVpF86+pXirzJ6RPYnZ3ZtiJnTEvnVNfRm8q4jN0wo/vopBiCxg3WAmeOOfN6P0Zr+Rr8z5TJe
lBu69O08JHkLdvO9uxkFCwFe5L4+wy3PFitNVabEy2QuNl6TaOnGrubDMSyS+8u9eChUS9TFlK0N
UFA0rOLZ+3/6U8CP4pg34Kr/++m7Wx4jhfEw6Q22x3qD4LlMlh+ys7Vz3+TMeFaJaTC2fgUfeAwZ
iDWlkBVOZ80JAIw44INIx+lgTGUHrKOxox7j1kz5Qc8xzIpfzJhGyqchDgCULErLdxJhnSuuts43
BYZD+inAXKKnevFFlMR4/9qu3dwWbnyNMQ/+0THxQVG4hF7ugMsh48fOVsR5G2+iDVjk8rTlw5tz
OOTAnatj2/T3/VZazb6sY7nwsOjon4Z8rSscKxKr/zt1i0ITMD8cCGME9ycqJQKpAOefE0JyQKZG
tvvExGlG48w0BFufSUwYhM741Q6p6Oh1ZgbDR2+oSFFHCeJaC8cZIi2hbix8cWzT6YYevreZ5N4Z
hxLZjDvD0iOFO7VezPsAnAXXDIBcSDanlmoZDe9MpfYrWKXG6fVkRWY0cMBxhr2lBJVCjsWm8uIR
cvthW6M0fAb3TgjB5oESieGmZPYwpCvwISVcSYfEtO1JWNnNJ1Hq9cGTSVGrQ8ArFHbxHyNiF7Gx
V98MLp2oEkndxuFWrlbOiLuXmm3T0Pwc4yNwJCzeIz+NCC62AQiaYCUT7F/iRPpUH0mxeIfdKJID
2NCmLZ9XdRPJfvox0KIFWpme0WW8hUliGLNNpZmw5UwZb7jrgDuDqg5sn+136MveHpfQBkv2qshK
uRPtwQ+oG2FPEeGjaW5lDp33XpEhD7yEWz386k++rw5Xp/ePuNDF4yoFjq6K/MaCmzwyYyCb6DY7
Ls0W4Qc2RW8dF/ZSuWOILVNLyIoNtkmw7vOzBJ4mjyE72npiS5ax6HRSTKZoGSVFINucYmnSfk54
4IFZOxC0ooBM4kLmeLuFqvUbJy0Dm3iltDH3wYuGM6XMbJ5oz1ztTCvlCMf5nCIiEIHdzvgYXBNN
MER5+KGs7o8WZnTAsqnSp6jMyPGPc5XStHtCx0O8+qL1P/DSgWVuec73iv4h+fw+iXsp46NwMcWP
DN8LMP6r5/U8BTfUr8LRcFD4DEtf7tAfgzVO51W4jLtPwq384pFbeHCGYQreW9FK90EaJB1nrShn
zW3VRGM3Dh2RS1eKWTb9x6W5k1drqB/zCU+dWgb1gEbHZ2hGDKPYujP2qMV1ytgBvFT0U/fl9+r0
mCBSabd2kunATaka/ofiHtT/5tUpA6Ds6m0eSQ+5JILE/MeFTYUEA85fJNUIIkv2mMQNyt+oqpYy
DK0lVYbHLH4iq2OQzzURn2ttDjvx29nEjoA0Lch2J2SOlsPKKFwtxj4RZIyEEF+NpKHU7EWVhzbj
bDZNPajqfowlY7odUJbMK/88FZTQ0FrOojJHsRHZ26bdp560QhK0tr1mJd4Hso3Q4UYyfwShkTLP
yrqzXW/yPjeMFB7AiMa3tfXImJGGk+cfvdWEoC2c5VbqaSFKeNdA1giCGF5rV5zax++0CUSnAgnG
f38OASs2kNnEZbzFezjFQU7w//dRctwtYFPyW9AowoSSbcxqgPuq5DFOpWf4uoChalXRTVoLXMGt
tzxqbmuVsYOzumzEPCqVPY3oZA61ANBGilrgIgi7FxyU5xMcTb8S3vfJgzJgL6v5EthStb5+J81k
5a2BUBOIjcdIBvt7qhE41AC6Kvl7698/zWMNV4JW9WiQBTB5c3/rxBU3015tXGgwqGZLaotXbwkN
pdStL9fVbqx/1IlhY+2FEUGnEGLzsaQolHj7Rl4UfNSoB7DIJenweFB0R2ja6C3c8+uQsHGC3eZm
vfh8/L9xe3Ky2NN4MMGsWOjiye6UVFoCbXAuUTuSGSl89+4GdtqnMK4hWMmqHL9cUQuQRUwG0usp
O+AMml6pmOsA2CwhH9i3aEK6Cmx3C+u4gfPAlVK+syrkr7aqr6eLzN5DhUGhlxh///QrscwRHS+R
QX5tE5wFP2Z90YsogCBjcGGQq4AIXqXAUVxNY3n03AelFf++axAIk+Z3x3roMvus+zwhfye76a1v
El8bFauTkqZFnfMOV5G5x88FXqrf6w79+yTUAKDnOBD9En/jFW5vFDVx/R9RUSRwAJLbIGGsCt7v
WQue3THVJK7lEY+54OAOFd4v3DpWUyuNvxnjVZqoKitIbGVUAzys+bPvrxNMoHWYMnXd/nOISzyg
kbAwEfa8EQdfCdAsppuHi1SlpEwdCs64fH2QjHFMZD8URKbUQ9dBIUa35XKoORPkEFjQVIzMEn9O
vqEq+85jvNhe9/jFWlbFmWBoU4XsWXbKGJlGPyZFt+49szV1b7efdqE3GktfP8ExksHwn5Ey0K41
wX+LGkdpc98boPgCKbAG1k5B7UCvNx3VHWgqWL+e3+OY34Bq1/xtX8aHqewgKf4GQc+or1Db2dj8
WuzainB+Ax+/tF9MV4ymLNctmsz0qLqt6h75ZcT7FYnzhECqdmCwbdaH14iQurelsRP663qGgRkh
rUcf4k82Gw4XnVssmJQfNK4d3DVQecxTOlqcoR37CIuOyWlYmDsK5LMpVyf0Py003xsjgFtwioOi
X76yh/fh1Luguf2ibpQr36y8aGQOlwS/HeZwXTAE6zvwiir2gGtQ/gpKwweQLzxh7gTrwbVHXfVb
L0uKqY9kVh8Zd7FIIdsoJFx1G4X22gE0s6vh1Bu4+gi8LSp4BnL11dI9XI8y773GnZ1dmN/CDZyX
Zdr99SYapmnzv2djqZ6s+VXxyWW1JjIElg+26ZxrHiAf1PtxiibWdfxfiNp/cvUkbCTZ+pA649/p
6QM2CzLDcwSfFrncT79fx7t3lcaaauFcH2NJXl7AK1hu4OlV+uaH02txStHmZlBppb8cP3lK6Pxk
hLMsdFfImb+uwCe7vL0tYk+JRDHED05br4UTLggoZUd7sNilszR9deOi9WopBCHCaT69kmJbvTaU
byG3f38nlwyD2Z1uxBmYI2Gbcaii2+zf9CTnd9rFjWBwq76KswOejsssCy1cUICbcurFe7QLXngk
rR889hkIcjP0eBT43nOqTd7l+4xq+59tiACZk91E6n8y2oxumdMmIem5mRyxY00HOb3YUXjH6tX9
jdjwyVVsYnz1TItUFgtzRIw9jlX+MUXC9nHCWKJYzLWX8E68Q4hQju+ZvVJsgV7YOmqSLEeXZCdV
6yZu/s1Zktrp+bUhZsxqF+2h0QWHRA3LaV7z5ZN5aateUQCzLYdgTe9EU79xrcHj8MRAkCaHh1I5
8VbEbFSDJJb3nOMOwDY8WjqkTmCsoQoYbGgTxdDeoes9rnwh9J7XIF4AuUV2M8yG+D4kv2x07fow
m71aYANhK7bQdq+yZ6HB8WI9kWiRGH/EJ3rQNqutTRzeDyZmKQgiBnmMp0n8S0uCdVSxScG3earh
l4NDv+bQVO2KWvcxdNZIbmyPgzTkzCeMkLlovOlR1HzjgZR+5E8iNSlooTsw7Y/5yKp1nROI3xsZ
Fy8yXTLWt44/Mho3gBaMfkgZIzfEGoeZv9y86jZyZwscY0A65wiRPqugPen7AizXifTRlE4Yf+QU
jrwBl/g6KioznTvle8MiMhCPKawRcGmrxRZoNheKky/gRQC3hE0hX11F6sYPjsNs/3rr0Z8YNl6l
rzbl2heFmKjDLQnbiRsx1KUJNxlAPYtGxdW8C8460P1w/U9ZC4K9zwej1kgCfnAoJgncV3vLjHv4
wE1n0dab0kxOzfjchlf2AdHchVW120cERI5DnN0gPevJe/UM+Yp5HvdXZFVmY3gXCMf4V2rE/Vc/
AH2T9Csctl5HuSS5Ui9H38PG5DY9xplnCVv8OzuEKTe2Gr4D8+ZpJ4lVfCgH3D2b2O5hBa4yan1y
Z2bb1ezkdZEqcwnEimSAJ3eAFo/c7oZU0jb3gjHi7oYkZRiYznR2W/4iV21FJ9TgaKvOqDctRb2v
anLZ+3p/euKnR9r7hYEmjnePA8MeV1tGw3g7Px/0eKZQQmO00O9ioDTg4o5YYLd/SUCrQtV29P0v
y7GswLqRqTGk2+0UMaB6s7hYP9fBOLNJwjDFAKq4X8j+yjK1ZxDDj7YG+kqQDITZOPXOLR9ea9yO
C8q5imlshVIdKeM6fvMwhZ7QlHiyDHoETAwTPNGGxPwZO+1Tggv3OcUm4DNf8/RFVXXNzzynPTuG
Oosj+/BD+2kKQUJ8WA/Zb4lKIweAcT+FmWPqJ4QSmcKdOkW67hdIfDvxnkmAIgo11GMeq/jJMtXD
ha9ZGgiG8t+ElcILTgGv8z2qVM3w02pGSONSd3szHcEC0NkT+EFmSfyog6uvTowFq8r5h6JVnNFB
r3o1SWBsiNfdF002TdTIbwawxXBiRzyuHr4t077ochGeUauSQi65xsHuWyn713d4tWXGoWNV+6E+
+Cw/2+mGhJgKr79HS2Zw0ld4GGeVbDyvONkjbYuSc0q4tJM33R+H0Ou9KVbpu/oHXPzjy6O0+2iL
cl0iWddWRppVXBny4AoOwB1drJzFWHkjp3pCJId7jWuTAXjiCNZHCiTZt8KEM1Df895xDoy5UGlZ
0skIZ5yUKP+L7FsaZF0dEZVV8y8hQTKYG83uhVgwnbxIwbqHq+yJq2O0/MEf6uqebulBthUaCuOT
/likiwQ9DIfIXlnCPQZp4I9zurCU0Cy/B9/ZXLJErn92T6zE1O1Dp5kyWh9BNYykxddj/MAKQdtc
ck+Br5VyE9Dfs8dDHZjNnsivQWGLcbV106mjA2RP0F7NanhJW9PXs2RskCWvjfGA8GjSKbHQbKMJ
NwKI+2Te8NEV77zqIX66VOyr9qpd7dvLhCrLMy8r6ZXAJiqL7Q6Gz2ld9/2mkFM+GXFWtYOIZEZg
flgsR3dXwUHeywVdvOXD0mpiK3/AIVpFv4w512z76uyeqsdbAMPnOZz8Kp1ve/xbWZS6HbRH6stV
+h2XMMYseUgGz3YKhHFe+1dEullgpzqLodSHG4g5fHdVSHKyJV0+Svcv7aAspVpfEM/ATqXsWJ2f
Iq5ZnqTiFK93XGICDV9vPTuuFZcbmsrCbNHOt3mlpE8QowzyfhF/Ouycd37pUU0UbR0Db5SgYqk8
0KxFN++HT1KpPO1dKytRCbAFWIJGa4Ct7B5/hcwd9o+La6e/tmEY0ZcZ1Ladmk5m3O6/udGtNlH5
VKTp5XHl2Z19oKQjyLk92sRtHBqQiCuU0cyt7xdylbTYXl5RM4+g0dgceJM5ZiCN7V9j/IZBWBZl
WMzm6XbA+NrMvoj+0DB2RHvRe0CbOiR11ktFbRE774yrI9LwJu7I29FSZ1bZ76knWvsaa99kvYBu
FY5XGzfbP4uO1VHe+8VMvwfwub5QCL2QgdyQmeFoo56z41dQxDe1VW6YATrxRMEBRLhQl9lI8uXp
k+k7edKokUA0FC6PzL4iocux8QoXrVYOWpEQb+RSO5cRLHcTjFCwPIQvHkKYoiHW1ZtnWs+rgJkJ
BiYugRYEPLcdwzGE+hROxZKiafJp5JyU/Q3tebI36OrmubDUcg3BfaIIisVGD4XlRSDOd4MkrrWn
CwBBLcgAAgW81wlEdzV/OeaQe05w88jHyHEMa38Nfr8JxS5DFfC4lf8+GPTa6abBrD4YQWA/it5F
4M8JcpY4NRyXoUMuDpQ8b/OwdB4a9aB0mNVfqsDUUozNtuCrQuwGxh8AwtSm5ni+wQib79cx2aCj
gABNIqMosTVKFm5O9BGSGOj+E/QIcHpquxK6nDnUKfVnCd+gkoyL+5Yg2CNLdjZJJ6kRsRxZUnmB
ZSCFriqTMbetv8etKyXyZgADS53o2lo/DUizXuxJ179HZMz/5Jag9tCSj5Yq8+g7CewxNgEr98MZ
uHZkIFpe+/gzJw/x2cMzRsjjIrhg2yxX6wgOdn+TLY50LC1o/vr2f1JL+iwgWP5lFZoEH1ph0zvC
wMkF6MyBeFZTyNokywjtfnNfA/j/PTzyk8QLjdAGNXsI6qUjzy9a0pzIIxzMDjmd4Q/lMABBD3bP
pLIoUaZRK0XQ4JUUCyzI4NYTvkC5RWyz9m0XFeYRBACd0oMhMk6Qmnpo85piFopdOWdB12394pI1
UWU5oNXp3VfLf34vt5MiwnBqjL2zLzgyt2FJ1UNRYZFNQxS9iST+gm2sFPtoeyfQAsDTPXoRmaHc
mf67qErnDRA6LRvpBDqeGluIegBoaKAz9NvqXU2TqL33/IXf0zJRyhJIHtkec1iCG7C6OQl5sgQq
FmhKIur85dr8tDMg9H4zRMSlvOx2jQbHW6M+MzewhXSuNfhe1p5PE+zp9pHrMI3cBSoffLSuNG8h
k2Vj1SsdwPZjrG9FFENqlAJ9hMYvRcx/qjdvmHE07eEDK/xZLnwKV1+EcaBvN0rImzIuoeMLzFLz
yeDaLyWdR7KanRW0fM3ok8I81FHclHljAnWqnq3tEZVVoEwWlIk7h6TBsTdXupbxBPmIwhQ4qzSw
cHeD4lTtWFV7UHZHGyKgH3GFfNHAGuypWQIACLoloAYpGxoR5+FR8y9QfvAxWjr3w5Nito/KUaAZ
ePHXFywtB5DwErni4dktpDbw3juQU2uOCbZmvXm9FhGXiYQdrCVP18EgPgeSTjU9dllrvOioSXPf
uKsDwmCwwGSreC5w2DDXpoZXGaEYm7GNnOqafXQP1TeQatJFnPttEkzXEdCcMwjJYjcBpT+Y4kPK
kIjXRJDzanb+TSBxCR8scX64bdLYvebC3Ek2GY9JoVPjeo6scguTrbPibK2iZfj59molsDVbS3KY
dAeTDpFU4hz3d7ni1Sl6vpzIzjdC5FSU23KOMrJHGvR3cwb9YXeGv4F/M1GKZcYv/MHHNYPsHP/t
UcvmnRZ0UOUsOAp984MQg4eyiJsYPWL879zw8zMqjUAwkqRJhOtfwXQNpzgwGsQ5CnRAWJJ/tSDy
z3MvM82jBOwequRIwoRikLjUGu7/RPKvmv4h9Vk7lvxrPRIuxMKC2htApgvEjzpX71megDCRIrps
w+hN3nsxh08gc4Ia1GQgaW5wlvbfAyOcRW4STg/JVNkl9f7gLu9fedf/9NH1hBxOwZ5m/BLQFKAe
eBlJx22LRvv+gfNO0hZGIkjqco7e5Penovh+RAQRp19kgWqJjSQHcSGJV1j1TRZhpKroV8/iHHZY
GyzxnlWJrtnuyyji9Ja/3hpaNy2Fec0gzzQJPaBO2AcicuY6L7rahGJ+6gQ+uPZTb2dG+ZaoZg5M
qYfxfwMINq8zhX48byXo9PsCiQY2eqb+QVq2nwGzOuQQUEtHMPrTKaJvpdacyLTxEZwx4DOz3JNr
X53LJTTbBTB8OpVFaIYZEhm6mFa7ct49zsHoPoCl9w6fmLVQPLcSw4tOCMnRP1Tpz/DH8/ReYesA
//aqfYZZrDrGppwsqXgXHz2te/8IYSSu9HjdEeAxGb0uKHFI2McOalo6FLkpBzTRXT+ogV7hHJGw
b3ZBUjwOA0t9KKQq4Kzc7YVpPypuWPqSjk2huJtO6WIMlQFvmw6sfIVP/0Q13pGl+ITf0M84tsIF
JIYjYW/po/60MlyfuMiCA+G1zfJ1RMrXZ2D5y5CXJ1PdaLtpvi1A2l35MqxZmtJIfQ4N+Z1jDW8s
QyfBl94XVscSqIihcKy5pqKEeOwWLg/HvY9efY3+6+eX43baZMPN6zHn3uaZM4GKqQzIo9ixFVL8
DoNFD2C84dxuQFFnNgr6SelCx+rr8biHmCV8AH5ua9dl66wNekQobf1JKpGk36aJlgjU1QZjMGZX
BuKiynZB/17tc6L8DCXHeqYrH6flvJOubmF/nM7FHW7RwHHyk4951Yny8w9qaJBklB+05912vsIM
loZnpv5WqTpPYxE12IuRd96W8Xb9GRIJYqBpJou5ax2rqFJ6mmIKlOYyPGg5t+4NyKuCNHt6zGDb
7BwTrbWLL3VgiwAn5BMmMqH0rd4j7ETolzZ2IP27qGba5xV6AgLspSwnGXzN4qrMzRRyG98PUXod
TjOYNH/RIpgNjqnILx/XeGLKCk6v+KgmvzA2YGgu+kl+MNzrtikwRy/JrKK0cEgey99CP6yLK1CA
ahbrVEroLo1eupr05uFkAQxIV68cpSkoMAoBI9GaP8YNMSkJ8axJUY90goZE2HgGCm82HhDJboOZ
hjjPMwV1D3jT6UNvFeg290xlVaippYZImYrTqPiLPnHAR3lV+RoupVMB6VCz8hQet5tjch9ZQT/y
d3KCnFleswpjDU5AXoySDMTjX2OqRCsDfY1Y6nlSPJZ68Ltd4mhiBoTt2lk9P0Lkf8K4WzHYmjLr
1j30+Zagk8ipTcirGFdVJki/75Ysz1l44WH81JCKS9FAjKKTVRsR8j+7Wqp9XpqiHPBCawu6xIz7
Qsv7TPs5qkjUN6qQiHueD8NKUc1ufx5BAKZblV/sOJqkFD5T1ASIRSJ9UOOkls6Gwg3KjToS55Pt
z0q+snpD8HLji7C8rKfQRYAzUwNfNMrjEr3MIZKjAZH6UZ3F/0rSkpaKt/lviNh/AWcJpzpWmp8j
74YELPlWOgdWT1XrA4tahmmyp/SnqasypVW5gFDEqlfYiNwodA8j3wQr3Dr7/eIf5UYoDN6pgcvd
oKiDmo4skzoTh6jXZ+td951uDkcQk0NsFSf5FKTUyh8zrnaBiBWjAIwJ5zgFn52tufzCtG3xOGxu
4QwZDTHWSM9+HdSash9iF8ZGvzwPkNO46Lob9/5oExqdu+q/18bLhUUpVzHXBYOkFOsLWQaFAzV1
DCx5VVxDMBkNmZ9X5VZmLcQ3CHjSxt3SUZzSAgY+O6wzgesQ+ie1HDl8hYd1E2aflpRa3O2IYlgg
8bLAl3Fv4IaCeCnLhJvoQxLf5WzwOhh1wjnYdqlMc344V4W/N2B71neDeEH/QgLkf7j26iDA6afl
yjpcKR5dq+gizCJQS0RBstqryihhj1wkg+tpY1LnHRpCw0NeBikanZ2M9R0rPkcc/wPpAcNgmXu9
xV8pjsaLq46T68DFr1tBcCpbbfj+EXFE2IYeCjSxdVUxEuvTRzsrmJvWrenMNNuDvZoRNze9feb4
ZALer/24ycXHOZpqNMJEbcO8/8Ziayc3mjSoETUAfHXdL1AktODrlYjhM51uTL9omKUzMtICZzIc
Fz2Ne5f56r9EN/ni0uz6UnMWipu0Yv3m9pws1le1onDM2rxdInkMCDBM1Dx6
`protect end_protected
