--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.9 Beta-4 Education
--Part Number: GW1NR-LV9QN88PC6/I5
--Device: GW1NR-9
--Device Version: C
--Created Time: Thu Dec 14 10:25:29 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity VZROM is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(13 downto 0)
    );
end VZROM;

architecture Behavioral of VZROM is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    dout(2) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    dout(3) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    dout(4) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    dout(5) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    dout(6) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    dout(7) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"9E2AC9857A68EAD3001FD1BD57A9D4A75B240075E080974B999B990B092B1923",
            INIT_RAM_01 => X"179AC0C6955DA9AB53165DA56082DD5F3FC55F63FFFF0560AE9E8C1EF4CD50AF",
            INIT_RAM_02 => X"28A87FDD5F827FAAD50023BBACC88A5240D3B18D0EEA417AAD439592C1C294E1",
            INIT_RAM_03 => X"AA89185FF3443FFFDD655A00FEE50A9753F9B5A5BDD602E6FC9C7C0B0CD0202A",
            INIT_RAM_04 => X"C1126C1D60EAF112103A3B2B9802006483726829C0F724E1127B817A1118157B",
            INIT_RAM_05 => X"581EE01464F32798B495246696057138F5A2F5DD4701B99429FABDA5883B8E15",
            INIT_RAM_06 => X"870060B279A696232CD54A8724925956924782AC0A713C1E10029538CF0700C1",
            INIT_RAM_07 => X"98B7DDE8B07DF7BF675000B8A6954CDF790187DB6753D19E77FD776898AD2D84",
            INIT_RAM_08 => X"BA88DFBF6EE2878FD294969FF6F79DF7DE6E4DF7E19DA397F4936D2EE9B51E22",
            INIT_RAM_09 => X"F2FBFFFBEF563EABFADBFBD8B613F71C2AD91A49D994B705ECFFF890CBA2BD5B",
            INIT_RAM_0A => X"FD164D880F09EABD3E02224D1B613506E3CE835D7EEAFF9C61CC4C795DFBAF7F",
            INIT_RAM_0B => X"D78BBDDE977A5F73A7D08E772CCF1E4BF883A8310BDF198530FF7772F8971AFE",
            INIT_RAM_0C => X"3EE80B453BDFDB19D527F9F5539328956AC7E5D0F1BE2996E33DDBFA355D13D0",
            INIT_RAM_0D => X"FBF6799FD00AF266BB975BAFBC572F17C5E387BB974E37F38DFCC197D8F312B4",
            INIT_RAM_0E => X"7CE75A9B9BDC91F93A443BB80942206E9640F1B4BE0BB3CB7B6DAF7DFB61FEDB",
            INIT_RAM_0F => X"40BCA00582FF6DC0678CDDB11F1BDA3775BBEC2493BFB5FEAF6C7B795FEB3BD5",
            INIT_RAM_10 => X"EFDC425BE002BC8FAEFA96F70F67484CAF3B804E1E10256CD28A262600008F14",
            INIT_RAM_11 => X"F3376A4873E4FF0A7EBC933B2D59EECDCEAC6E4F339AA96A7B5CC69DFC1D27B4",
            INIT_RAM_12 => X"7BEB5CFF3DD975ECBFBF6E3D1A83818926314B174348F7BBE1D0FE2C9FFD141E",
            INIT_RAM_13 => X"03EEF6F50A502001C20210088086038003E7F50EEF7B4EB7AF7587777CEE6AFF",
            INIT_RAM_14 => X"F299BEBDFE62276EDFBDEB7F3623C00280D2DDFEFDE0B88DDAF7C9BB4FBAF7D9",
            INIT_RAM_15 => X"26AA686F9FA7A524E7DDFDE6CC2C79F3FCFDDF7FED3DFEFFCAE4662E3C78C677",
            INIT_RAM_16 => X"211092115827B504106A5DEAE29F59569B2688135B91155195BBBA8EF57DBE88",
            INIT_RAM_17 => X"22222224924F14F9C19269692B548E9098204960DD8B5DAD1058C64E24022222",
            INIT_RAM_18 => X"2247C2DCA4ECC89703C78A224F40BA5D2BEEEEE7D919BF1D4F2CFF9931843D0A",
            INIT_RAM_19 => X"C036D2FDE0705521007A28009201C20401C596298FB5399D2A5C6C224D00B612",
            INIT_RAM_1A => X"A877F3BDD6FD5FEB79B1EBCA3BC209AAB8F80FC894F2BD3C143803EC5F6436E3",
            INIT_RAM_1B => X"AEE8822485450EB1B4B563FE9F18F497090C69C50BD51C2D5AD50FCAB5E91CBC",
            INIT_RAM_1C => X"41BFB2FC1D8FC0F1FF23B7C1E6B8ABAA748AC8402E350A0BFD6C4E4ABD406D54",
            INIT_RAM_1D => X"FD6161222DF41471A98EA9406EA3A4AA01D4CD186FA7A6E158BB03137ABFFF7A",
            INIT_RAM_1E => X"8AA8C21B28D371E7D1FC5FF78CCA93AB38E4FDB74E44517C84379E5C78F3D926",
            INIT_RAM_1F => X"715F2B2F920421424048C1C7EABE108AD68F8FFDFD5582178B77FD774288A836",
            INIT_RAM_20 => X"9AE3420150428DDF3F94385618293144C1E2B114AFB8DBC20EE280B89176E9A1",
            INIT_RAM_21 => X"6912C4ECFE791E5031751A15461DC2B435D1007348C4B08FFBD00047115347ED",
            INIT_RAM_22 => X"2AD6BE3BFFF1BA3AA45C62B053D568FD17CC03BE2D0BFF3B847BB9D9FB428403",
            INIT_RAM_23 => X"DBA70BEE56BA27D56BDCEBA875FA93613B2A412A34D50293F4AF021A8D5BD7B8",
            INIT_RAM_24 => X"645ED86461D894240802A310976FB77BB9EED05BD670DDF76BF56302010200EB",
            INIT_RAM_25 => X"F386EFDE857B7743E6BB334356F57D4ED68E9DFA5E5F3DDBFD5BF9611A84B1A9",
            INIT_RAM_26 => X"0BF7E3EA779FFBF254BFD79FBE5FA9C0D556AB140453BE68000448EE77CC2B5C",
            INIT_RAM_27 => X"CF067106D9AF575F321957BBD566FF0C956EDDDE3C63FB9E9984158314B59456",
            INIT_RAM_28 => X"7AB890AF87C5EC469D52B5E854F56533F0109A3BEDF72AF5D7E8D1ECBB1CAA77",
            INIT_RAM_29 => X"3558E86BF898AACFED8FDB83A37DBAF45A353FF5F512AF98F115DB6B27CBAD54",
            INIT_RAM_2A => X"6D63FC7FDB675C7BA1BFAD5116366ECD0BDC83765C16FDDEFF759C774A1EEFED",
            INIT_RAM_2B => X"00B55C59BE3D5F4EC35663D20F2667596D41EAD9C78FD7F5563EC5E3FCA176FE",
            INIT_RAM_2C => X"76215115061E41B9B6BB4E9B24C92B5FF098337AFFF573747DDF1FD5FF23C035",
            INIT_RAM_2D => X"CD654FF8A17BA057FE78208585AE12457CAAC108020A892605000282C5342AFD",
            INIT_RAM_2E => X"1DBC042DAFE69767BF9E0D751E5C4C29021069AFABF72B5D17133B9FB7AFF0BA",
            INIT_RAM_2F => X"4088260024F215B16D4E53E049AB5349A3C1CFC480B376CCCBD40188090276C4",
            INIT_RAM_30 => X"377A6ACC0460263195045E724855AFFA49084043262A6E3B92421A4AEE0022CD",
            INIT_RAM_31 => X"0B032ABCFE6B6AC04FA149021215240B4A484290B7D0CA79FA15B184A38123EA",
            INIT_RAM_32 => X"1B05E8E3B47A15611C09B019C90620D802097601825C6C00C313547BB32E09E3",
            INIT_RAM_33 => X"5A4D497E2A38AD7FFF9A38820FEE7A4B47FD3CBC7E3FFFE4A31A0FDB28E768E0",
            INIT_RAM_34 => X"E493E278FA9EF7E1CCEC53702A80045E784F131BAC9352239F6BFD2D1068BEC9",
            INIT_RAM_35 => X"7AEE60D30A908721569109A0D340CDE703F0F287958080082110179B66CFEF3D",
            INIT_RAM_36 => X"68F7F359970FC10756BF1F3979AE79E2E480F4FDD5F7899269E4F847B7C01B84",
            INIT_RAM_37 => X"4A8AB0B0635F5802C580B0638CC7FA2B8E6556EBAB9FBB3DD775D8875172FECD",
            INIT_RAM_38 => X"F85BC642D0A168D421FF44341F467373737F7756194AB55C4FAE3C6E1E832A82",
            INIT_RAM_39 => X"F9697FC800189055AFAF5E424C807E63468DB8F087F9C9A90EACA3D019AF8DAF",
            INIT_RAM_3A => X"B1DD359ACB076EDE0C6EC9AD0E5027B7EFDDA3F3514324460034065DFD918F2F",
            INIT_RAM_3B => X"C08C2308B9DE71E2E080108C371DD7C07A7D77AC53FB9FF1B268D170AA548B94",
            INIT_RAM_3C => X"346628D6AB38F3E7CFE3104417FC771FFFFFFEBB7CF7F1AD77FDEE3F881CE739",
            INIT_RAM_3D => X"557E48B37DF232D3B2D5329E935F5347348F593A2D91D4A6F278B66AA26F3329",
            INIT_RAM_3E => X"022491E299FB47022DA088368CDA32BC444198751D95DD16817F94A49CFBA944",
            INIT_RAM_3F => X"FFFF0000000000000070801A25CD128057BDB691FE7F3D1AC68C4B906D516082"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"084738CFEF89F8CB0003043ADFD21DB81214E311121915C585838191B39301A7",
            INIT_RAM_01 => X"091900B66C77F23C83243194B9C5D4C39FDE77AFF20FEC5D892DA1D53688BBC9",
            INIT_RAM_02 => X"0A022A08A87FFFAAD50054A8AB449F9A00813B8BB04E006063C3031301B5E14F",
            INIT_RAM_03 => X"4F9091C00CB6680011E636C5821599E38952D9C6207E290082A4882C3412682A",
            INIT_RAM_04 => X"CDB9EEDD76C607394B9CFAC6037659A265014142991000ED54484700637B3F02",
            INIT_RAM_05 => X"F98BB6D5CC03C8511902D5AB5A37432713656C008F6799A1BE81894C14AA8933",
            INIT_RAM_06 => X"C4802210092DC022135DEEFB820809E0218A9B397E3A64B35964FF1DF92C5D9D",
            INIT_RAM_07 => X"70B7F8D172A6D7C2FFBC4033E41608BB831525DAFFDB3DFA8650822832929424",
            INIT_RAM_08 => X"0B19CDFFC186A01F8E738360002C0DFE68A68E0080360841180524430108F14C",
            INIT_RAM_09 => X"2927EFFD07DC43FC2C34AD3809FFE16BB87B5011ED3C1BF4BD50D1ACD0A7C7F8",
            INIT_RAM_0A => X"FB5E9644E9531F0965EA4801E5D25A719E27F729C11D2431B21DD54E28046041",
            INIT_RAM_0B => X"0073A83553BA071145A6016821802A1D21719EF3B0697458C4BCB85399963B48",
            INIT_RAM_0C => X"E82CA1E8AF4031D69C580B42E9DD4C38ED582F440F97E8CD9D33061891C062C4",
            INIT_RAM_0D => X"24082769000023100B33F4401E8A07A1B0B0481DA387F841FE11F4987B025704",
            INIT_RAM_0E => X"05B5FE96024099796B22DC68F6FD1BDCF9F0BC9C27EF01B825E0248626370955",
            INIT_RAM_0F => X"CB1815B79610D8F22E47105F7E7E002C0262158018707C8020D9900048109032",
            INIT_RAM_10 => X"A6DC8B322634E9A442F4699CD42F7B6A77E839E061F13C8D24126E6EC4444864",
            INIT_RAM_11 => X"D0B1111C6C0C36BB2123268345C4D3E21136C8C2FAB4EC934C83736383641C41",
            INIT_RAM_12 => X"9D06400084A0061386A501E742F0934D72C052A929078C81964A457A6094E9F4",
            INIT_RAM_13 => X"201210284A483020038A140031A54E800EFE6A0321056CCF788C4F1238F7FB20",
            INIT_RAM_14 => X"5780BA233405EC31100230484003F96F88E002C0341D852B00802C4D208158B7",
            INIT_RAM_15 => X"AA445B7124880256040810B8CAF41B49924471162040D0655A0C9CC0DC9199FF",
            INIT_RAM_16 => X"00000000080B2B000015D9A29C6ED6B604080401497AEBE7FB050450403B9D0E",
            INIT_RAM_17 => X"0000000000044978CE8432E75D170300280000C06892ACB100108EA60A000000",
            INIT_RAM_18 => X"AACC7ED8263EFF1FCBF00D67423CEC450514142FBEF873E0F99B50050148B8AC",
            INIT_RAM_19 => X"001BA01B88A173076DEE416D25B64EC0C4476891BA005DC79C13024797002566",
            INIT_RAM_1A => X"F9E2083FDFF1202508936634C80F3E73F150C6010E668671D2F0DA000CE178AC",
            INIT_RAM_1B => X"C18D1BF7937DBEF379D9878CC33922C8659DEA3727C8212F9FDE157B73003CFD",
            INIT_RAM_1C => X"2E014948C7133FB6C2640B0ACFD27FB01583D4D9BC37CEB629273F29EC73FF73",
            INIT_RAM_1D => X"07ACDA3BC066C806CC32082062E6294CAFB95FB516DECAB7F7EE726326CE0289",
            INIT_RAM_1E => X"598B35259E9356D9361628AD1B817B13D44D06E044CFB5AE74D3221A93E8A25B",
            INIT_RAM_1F => X"EF4AC6BF9ADDB2EC7B1D4713678ED69D18F330A1424C9A7C461D95D86BB8E2CD",
            INIT_RAM_20 => X"58CB949723619204ACB94D395961A7C83F0532926C5FC08C3DCC4F2F5367A27C",
            INIT_RAM_21 => X"8D7B0D7B609A655864F1E84EA0D03E4D932302699ADCDF94BF5113DB5964CA46",
            INIT_RAM_22 => X"BC3FFC844C8FCC45382CEFEFFB03C4496A3D80FB4ED63DD0B9F10AF66DBE7DCD",
            INIT_RAM_23 => X"36002018784E49EBBC559F5F8715BD8C4FBB27725FB72CDA49B2DB263884F9DE",
            INIT_RAM_24 => X"9B931889B643D9CEF7DC4CAD9C1A89960010296078D2B009860B8A3FB52B1120",
            INIT_RAM_25 => X"AADB18EF17C76DB87233C336F90FA3A123941CA7192B453411E4C79FA57BEA5E",
            INIT_RAM_26 => X"3AC86C114E299F6AD8400F32154122F5CD62E43AECDD40F40023B10C8772F65A",
            INIT_RAM_27 => X"3F6F672910951A71E821C0D6FBE3F99EB227065525C75A3DB67D9FD29CF3599B",
            INIT_RAM_28 => X"5B81064178DDBDC9D4E8085E9D2796A4E316BCE7C90A5C9B211E16118C72CC02",
            INIT_RAM_29 => X"BF634BC2261E3F8B1290A26C5952188190EF0000E163F959C6362DE68E8FEDCB",
            INIT_RAM_2A => X"F54717A184B9FDCB664988EE6E4C51505E1124FD4C82A358AE5194E4BFF23D21",
            INIT_RAM_2B => X"FD821F3C21E84127E5F2F9710F3AF361AE728F638CD7792A78E20AFE68B31B9A",
            INIT_RAM_2C => X"8D27BE0FE974587C8A2D786CDB36CFB7DB3418054E6FC117002C663B3E3C7FF1",
            INIT_RAM_2D => X"272BD0AD3672CFA4300D6E6416E856D612F0A7EB933E2D725DC6244FCED75F3E",
            INIT_RAM_2E => X"264692819200B093000DDF6FE41E00BDB35BE58A3DE1BD6638A8444C085214CD",
            INIT_RAM_2F => X"99B97B6CCC192A67EDD0F07CC5B324C5B60B1FDD6EDBA74E90C5EA39FD661E4D",
            INIT_RAM_30 => X"408DAF19D6DECD7B5E2BC23C217DB24C92D6936CC752FA4EF1C959240B6CCFD9",
            INIT_RAM_31 => X"602F6E5C9E66664982ACC73FAF7E5EF7E4BDBFFA4E53EA6AE13123B04FB2931F",
            INIT_RAM_32 => X"5838BB8428F363067D91E578F420E4111843044A90C1C8F5487B299897607907",
            INIT_RAM_33 => X"8005863B3AE162CAAFC47B89E415886C2122905D88D99983CFA917A8BB8851EE",
            INIT_RAM_34 => X"0AC4388101A05405245386EDDE5696C221C42C08B020F1968EE86CF07B66298D",
            INIT_RAM_35 => X"6ECD6644F46BCAC5F6D2E7B39F6F1039E8020D10384964EE92C9D8048550A142",
            INIT_RAM_36 => X"03C208C5B02818F4CD52A91AEF90D650805F5100BC06EE61A276E7BC9C7B2E09",
            INIT_RAM_37 => X"9092B2B365B95970C99BB36504CE079C2C82AEA2988DA867B0EC3BCAF3556ACE",
            INIT_RAM_38 => X"007AA28BDF45ECC5B7FFBBF064949545454554622CF311852F3724CBE093BC9B",
            INIT_RAM_39 => X"FE56CFD28B080D98F2ACE110333FC1BD9B7681472C15264E6F96B23A87B4D75B",
            INIT_RAM_3A => X"445DB365EFB6B8D562C83231F527CB4952A375AD9F947ECCC9E6F8ED2B133AD1",
            INIT_RAM_3B => X"DB739CE7309EB5F6E77BCE73AAE00C2FA881E33F8F028E638721C346F379934E",
            INIT_RAM_3C => X"5E2213FB8FB76FFBCE5CE77BD373B2E7FFFFDAF7BCE98B2D77FFC6FEEBDCC739",
            INIT_RAM_3D => X"A5B095110A2B7341B03F3354B14402821A5A86211E8A04C9863B66CD06371164",
            INIT_RAM_3E => X"6649B279826D49665BA79977EDDFB981CCF1DDBE7D6332A7349FB6782D1B0022",
            INIT_RAM_3F => X"FFFF00000000000000124A3931DFC048CD21C75224E271272893BFB37D920995"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"76030E4F8B41F32380058003C046930A5218350037281206141212B89A9800C2",
            INIT_RAM_01 => X"0026C1A27618CE240547193471259A800A9756AAA8078BF16D2C6D40BE6EEB6D",
            INIT_RAM_02 => X"02228080AA2A7FAAD5003E99B054074800063C890D120187FD7283A4C12372FC",
            INIT_RAM_03 => X"EA18C88046D0357C08317C4DF1F42A956D9CE1F81B7C0A007C451CB00C10A02A",
            INIT_RAM_04 => X"4B29209104A4223E63A04389E67211626471006A9187142976438200115AAA11",
            INIT_RAM_05 => X"618B223468091E438FF6607DCF6259287496181847453CA12A2109680C19C505",
            INIT_RAM_06 => X"0380030024990B61A50CE650E38E1466A109122C5433390A1040AA19CE421111",
            INIT_RAM_07 => X"40B6D9D912ADB7D2AA8555536D068EDB2515C596AAD2B2DF0F5C8CDC54898824",
            INIT_RAM_08 => X"502ACDB7708AA7AF04A16F0C31A03DB64046EA31C00469815C0BAC33EA2A9628",
            INIT_RAM_09 => X"2827E9FC0952C15400024202C251ED6149CA5415E1515F14E45658A8D5A757C1",
            INIT_RAM_0A => X"F8559483485D8D0D369206012032B0A0932824211D2914082C11110B2074A244",
            INIT_RAM_0B => X"7F8F531A337C2F8390C4043A82D520D5B90136D9345A4C1A6486534415BF2F6E",
            INIT_RAM_0C => X"BD64A26AA3EBEB2D74954A72AA1A7C52AD5A0D9740DE37A0E121B302E361C844",
            INIT_RAM_0D => X"A00BB14568028944B7B665262EC80BB5B1114C2DAB88BA422E91493A63569345",
            INIT_RAM_0E => X"FD6165B18A30B4D3A176F6DDE73BBDC867889BB17E2C6218090A2E2EB389A812",
            INIT_RAM_0F => X"C30C2C05850FC322EADC9AE5762C3672CF9A9E7317403683386DF28E7F5CF808",
            INIT_RAM_10 => X"0414997AC33209079B99C304380A11FE937871994CBCA03DE400D848EC6CE824",
            INIT_RAM_11 => X"870184DAEB05D6EBE86F227A1803E4D88E44415E1EA13364682F0C66E04A86D1",
            INIT_RAM_12 => X"3119DE2B20716FE541F69E32D03291E794941A42A63287A348A9C0AEAA520A1E",
            INIT_RAM_13 => X"D184218012482021800514182003CCC00CB2740268015BC0D738D800DC33373F",
            INIT_RAM_14 => X"05081631C773363C9FA2566F8C03E247B88161B06C85214C06C392019C3C7B91",
            INIT_RAM_15 => X"DAB9D6225984128962B33B2EABEC148571DDD7750B2381D9984936092352073B",
            INIT_RAM_16 => X"00000000381EFC000013715B6B976ADFEAE96C00B69F01544111442EE89DD409",
            INIT_RAM_17 => X"0000000000036B11F80406DDDA6FB5006800002064C7E2C600273D8A18800000",
            INIT_RAM_18 => X"AEBFCD2F39FBD642236758A170B84761011045336EE93BE8A98D012DDD3F02D7",
            INIT_RAM_19 => X"80E7BC5E68184570480012032C81260E2C6FF8A81970500A9484544246800346",
            INIT_RAM_1A => X"4205B624100A07014764EBC2832C358E081026620615717C1030430432FFB8C2",
            INIT_RAM_1B => X"FBB39C798DCE309185396B9210001405410C46144145452E9D0BA85E67888261",
            INIT_RAM_1C => X"3C1991B3C1E9D2E179408D56A149002D4243A41CC2C2651C0026326C907E9E33",
            INIT_RAM_1D => X"018103A0809491F0C121B5004888EC6626681D71743F3E80A54A315654BF9B33",
            INIT_RAM_1E => X"0AB00D07860D91F6A18A62D00080168AE20D00A34213846A75C4211AF3EABAC9",
            INIT_RAM_1F => X"F93DAB405801270B70880EC4C7621004042FB04C9A448AAA0928F93F4310E28B",
            INIT_RAM_20 => X"D60652D54700A0DF3648EBD87248E58062448486EF74C756F60014CAC4C1E819",
            INIT_RAM_21 => X"F85ADEB6186B301051A53242E49806053D3504225C5004A33C999950401C5149",
            INIT_RAM_22 => X"A26940722B117609AE10C143A3DDC2C1ABE50022EB68B2016CF37D6C138E155E",
            INIT_RAM_23 => X"0B9B624F61903B2ED502F4B575015AA408AB62A214B26C072D27BA0800412C09",
            INIT_RAM_24 => X"866BDC9C62588AF299EEE7C186CD801B6904034768F00B1119428AC94D8A102D",
            INIT_RAM_25 => X"C75E0EAD9483F651F318B520A9EAB2A70DBBC340F72F470F0C1CBDAD691AE2BC",
            INIT_RAM_26 => X"7D0FCA0146418002808E50BC9966633840C20358F55042F40076E1ECF75EBCD1",
            INIT_RAM_27 => X"475AD40CD025D601296D1C3B2AE00088A4E0D180050030343A0D0A588CA44503",
            INIT_RAM_28 => X"5028842308153D0583936586851481821582EE40618F34EC17C661398E416A3E",
            INIT_RAM_29 => X"2A026A88C180F5141B2B331E36E1800560DA638141595D10060294488E644800",
            INIT_RAM_2A => X"9C29849107CBAC6267817CF9982699CE551D07D6155AD88ECBEDA136951E3DE0",
            INIT_RAM_2B => X"1160100031373C62A27539EFF01C346D61736993D304AEB0281C9251B9A4D0EE",
            INIT_RAM_2C => X"B8476B4A8E59500B21F32E1C24892D97B8B863150E1280B04C6860693D23A32F",
            INIT_RAM_2D => X"692A9E2B9563EA231E1B6EE59818C493F65B26EA3136BA7E784366CD4BB39779",
            INIT_RAM_2E => X"07F680A10C1461FEBF1046862404040C20430969A6005B19B81343370B506703",
            INIT_RAM_2F => X"15087A2228190841A902A06E8522508106109A9F4652D58AB317EA28F10436CD",
            INIT_RAM_30 => X"10F62A59708AB410150A820E001D087C51CE5228C5309B6AA100502C6A620351",
            INIT_RAM_31 => X"B00B4E316A43448D0BA884235AC214AC64294852D5D2E94AB92510582BA13ACA",
            INIT_RAM_32 => X"525DBA35247B42415D04A5583800A008EC02020D80814426C05A550C654220C0",
            INIT_RAM_33 => X"50058F7B32884A4006CA3A81492E930A4125083D308C6C62A93186A7BA2A48EA",
            INIT_RAM_34 => X"AC9742EDD83B7768480554C80A1180D008010A0583A1A9B4028812A05244A2A1",
            INIT_RAM_35 => X"7E8F40F04A52C220641445091B4691454350DF86BF586C6090C8C01B6ADE0BEB",
            INIT_RAM_36 => X"00C5B680214C1483847E3E035902B1C22C48FC5F2851A90638D2FA0737DF3B89",
            INIT_RAM_37 => X"D0AAA1A1410D105881092041408680202EE27CC3D0003C7B21C872C2D4602A2D",
            INIT_RAM_38 => X"3C309080844042BCB555E32CE6D6D7777777776B7D4B5DA6A2B02EEB10A03EA1",
            INIT_RAM_39 => X"53611A9ACA080CC81006B65004A9407385CE4CDCAFC549E14B1ED55A8508850A",
            INIT_RAM_3A => X"0155251D7217D0848C680A35AD32AE66AD5A4103A5A6B4EE8CA34571009BAC2B",
            INIT_RAM_3B => X"DBF39CE7295ED5F6EF7BCEF39CA0DF247E2F5C695452366A244D1244A452A846",
            INIT_RAM_3C => X"C6EAB4A7BACBDC1DFE5CEBFA150DF66BFFFFDC6FDEEA9A8577FEAAFDEDEB7739",
            INIT_RAM_3D => X"958731F575D3E71B39DFBB2837294D2BD418A0768127E9FCF6FEFCD756EB7578",
            INIT_RAM_3E => X"460930B10A1D4546122248C0CB0329088CF5574621C4E3352506B6A4677055A9",
            INIT_RAM_3F => X"FFFF00000000000000040232005D8000443ACB51004021130A8912B109900984"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"1F337CC9F1D55D60400FE6840024A21444883E3323EDC60EE67666C644C41412",
            INIT_RAM_01 => X"09E1C1E9A1DADF6668ABD2639D44A8F4BD6EA006F3FBCFD9F92A6D08DF096935",
            INIT_RAM_02 => X"88280028202A6C6C6C6C53472086C8400040BAB975F400F647A58363C1E22721",
            INIT_RAM_03 => X"C598CDF452D9644A1F7EFCDD89BBEA878E1F01FF35D5B780C0ABDAC1886BC8A2",
            INIT_RAM_04 => X"6DF3C01E00F392915B4045D00375C44174C1B5121D0C0A0E730635CD1A9DD5C3",
            INIT_RAM_05 => X"7AE6EFBB97488118AD97AD45E67EB7FBEE8497166B0A6C389F4CEA576BBB85AD",
            INIT_RAM_06 => X"0100623254D362ED7DCCA67D20820406880765C9AFA2EEDEEFAF17D5BBB66CE6",
            INIT_RAM_07 => X"A0DF7FE54C7BE6E79ACC51991A61335CD91B32A79B95A4044139977CAB6D68A0",
            INIT_RAM_08 => X"88E73A68F818B66BA73D97F4BAEA37DFEEAB930C109DAEA1C4068AA0800CEAC0",
            INIT_RAM_09 => X"464F91A660BD2446729B94BF6CACB672F280182D76A0844BC21BBD1399D57780",
            INIT_RAM_0A => X"54ECBD87A617D09EFF79CE0731F3435D778718F3EB57598CFF0DDDBDF3AD5EA2",
            INIT_RAM_0B => X"4A777D3DBE95EAD2E775438EC6D772AFF3F088F3B915BD7CFD6B65B5C4697DFD",
            INIT_RAM_0C => X"1710DA9E95B2EA5D73AFC0E6C3A4D8ACD71ED7C76E779F71DCC3D714EBA1B3F4",
            INIT_RAM_0D => X"CC4E5EF64006CC05B56887FBA3E46DE95CD87187D9E8EE9A3BA49406B995E89B",
            INIT_RAM_0E => X"83CA27AD44E2F9514FEFC670D6BD5BF5EBFCB7605097F9913A049BBB97D3F37F",
            INIT_RAM_0F => X"7A8C24BE70396DCC738FAC6701705BDB5FDFBCE04EC12BBEBAE08D8E80DD8632",
            INIT_RAM_10 => X"32C4AFE22EB958152F5A260D53202A5C214DBDCF08291021326A2524FD75507A",
            INIT_RAM_11 => X"920B8052EC0F129A101526E22A818CCDAC8748F251800168C4145F29E1385D19",
            INIT_RAM_12 => X"312FB3B820D5C40747DAB88A9D298F22AC198D0E1E8346E5CBA7E04D4B600D04",
            INIT_RAM_13 => X"1E95A2D04400204003820A20E123078007B3710848123AAC182A288344F9AA70",
            INIT_RAM_14 => X"FC848D539E45DF8AA8615ABC9403FB358B20D5215A50B3B72B4E5311B8A0F46E",
            INIT_RAM_15 => X"EBECDADD30161B69B0DD0D7214543A10D42B0A512DA5CAB40A875FA0815FF80A",
            INIT_RAM_16 => X"00000000080A38000028751248044194430C14008012EBEABBBEAFB507432B0F",
            INIT_RAM_17 => X"00000000000449926806039D5F074B803800000030A080C2000E6CC60C800000",
            INIT_RAM_18 => X"CE260C2CA1689395741D55667F4DBE6C2EBFAFFFA7A7AEE9A958246C32824205",
            INIT_RAM_19 => X"80AF5CEC872D98DFD76DE6D524CF057B5E9F2E77D8EE5B50961060621F809674",
            INIT_RAM_1A => X"6D9FDE83EC01CA9C8AFD1A6B0AEDBF5D4921271DE415E37AEB303DCC76CA795D",
            INIT_RAM_1B => X"989F5F7D5EABBF794D7F9AB724DD7DBD9646612DB827ACBCD933519B7BB0C662",
            INIT_RAM_1C => X"3E03D7CBC3E0A56A55FB1573396983DA0A3D6A1B47E0AD267A9CB47F49D6346B",
            INIT_RAM_1D => X"9DF2EADD21B9674A924725C09FB7EECFAE8E4A74B27F7B792E51FD90C1C22FA7",
            INIT_RAM_1E => X"671445DB27DB9ABC2A2AEB7C4ED7EED1B5647D7807FFCD5F79D491A1EB253E49",
            INIT_RAM_1F => X"DE79FE500B3F8E2FB6D62FDFD5FBEBCE5F7E3956EB7CDB4965E04757B25758CB",
            INIT_RAM_20 => X"EE9CDEAAFAFB7BEF42FBC7FB6E7CE9643367ACE055352AFFF3112773BBEBD28B",
            INIT_RAM_21 => X"7AD7355755DD24E8239ECE717F6A5DE3B1FD0E08D66BCF7AFBB817BA7FBD3DEB",
            INIT_RAM_22 => X"FA8843EAE65645BAE411BA552151A152074B8092D6701057D288EAAE57D5C3BC",
            INIT_RAM_23 => X"A040351DC2D5C08087200446FE853C0BDC79DA9DAB328563A8EDBFDCCF470892",
            INIT_RAM_24 => X"DFB6F0D793374D4F53FFC7F74F5E623FA6178DCECA4BBD333FA8E655963FFC94",
            INIT_RAM_25 => X"B6891D103E11FEE7E39CE79A2B82DCD12B79AF9772B22893BABB945FAF2D5FD6",
            INIT_RAM_26 => X"F64A1D4C2491480A7594B81050C0782F1CFBFCD743B7306200AA05F7EBBDA0ED",
            INIT_RAM_27 => X"F3B1DBB7C8F873BA169BD5EA08C83FF29DDE57002B98B012248B8271CBFFFB27",
            INIT_RAM_28 => X"9DC50951BAA36EE923BCBEA6A65CCACF9D2D6C3013DEE5CB7BE22A8CC1F75D0D",
            INIT_RAM_29 => X"3DB48DE376E3E520ADD775B95A6A6A1EDA6DA4044DB44B7FB2D357FE67C45FFE",
            INIT_RAM_2A => X"3AB3E9C3C5852BB56363FBEE5F4F3BFD20395CDFD2BB62BD19DF42FAE5E95696",
            INIT_RAM_2B => X"99FD51F65DA471543C4711550FBD18CA93BBB7B3F4760BFE892AB3BA93C9EBC5",
            INIT_RAM_2C => X"E846AAF2E1D5BF7D73EABEFCFFFFFCD357E73F4886EEC36FC5183C0D1B5537DF",
            INIT_RAM_2D => X"D8E490937D95E7680880CDAB2EC12497215526D1B5F532385A76A75DBFCB55DB",
            INIT_RAM_2E => X"B77AD890FE04DCFFF0676332BD3302639EB99AFEDE14B4BA22FE5452CE54E787",
            INIT_RAM_2F => X"E8EE2EFBDF54FD3D47A97D4CF4F9FA74F2A4A54C557DBB5782D49ECE2AFB83AC",
            INIT_RAM_30 => X"004517DDD2D94D0A4E09F06E04C3F42A79CA531A1F3BC9007D2C4FBCD7BBFB8E",
            INIT_RAM_31 => X"38B2442EC3BC15CECB42F6A739CEF395F5E779CFC9E548B311AE181C31DAB4FB",
            INIT_RAM_32 => X"67D7BD87A6B7AAF18EDC4491B883304C0F41D32DD0766636E898C6A46238B5B0",
            INIT_RAM_33 => X"5007CD5BF7455F9FFBA35D69BC09074AD521142EC904445355B9DA26FD8F4D77",
            INIT_RAM_34 => X"2CFE5FCF9FF332767CD3B59C9B1DCCDA64CC8D9B798051739AE692D892C6A121",
            INIT_RAM_35 => X"B1563799926CE2331FCF85056B9F8C5CBE679C3CB3D4AA1DA9543C1264B1A30B",
            INIT_RAM_36 => X"34DFDE761CB778D7F064323751F1A51F362D26133728374B0E0109210918A48C",
            INIT_RAM_37 => X"407C9B1B369E6D6F6CD81B360F6A4DF0B70515455E9855CD3C4704E20EBD3112",
            INIT_RAM_38 => X"773F36E67E733E7FD8AA77DDF2D26E9F9E93393329419CD052D02ADAA47C5E79",
            INIT_RAM_39 => X"FB278FDA298C2EEB1FF88DD027F261FFDD3F8583E434FFE70EEC8DC88DF39C16",
            INIT_RAM_3A => X"C7EB9EFE5575D0593B9B7841D0BB4F7BF56DB36FC9D71DACA923B650FA8B24F1",
            INIT_RAM_3B => X"DB8C1D07195EE5F60F420EF01CA99986930B6CEFB49E9AEDF3FEF9DA71387971",
            INIT_RAM_3C => X"64345C2E30FDBFFECFC31DC1F6FEF6ADFC19002FDF7771AFF7F06EFBEEF7B555",
            INIT_RAM_3D => X"84CD191A2083612B3153B180118B1048F29D50182002800AD22C24E402221A42",
            INIT_RAM_3E => X"05ED2E25E048BA05ED1F27509D027CE4A24C9D8522E823ABC75A22A1357280C0",
            INIT_RAM_3F => X"FFFF000000000000002DB12F431A819FB808820E93A994EA4077712E868E2172"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"493AFF1C9BBB9B4B40027CC36A74615C86A0B256B67CD002EA7C7CC444440445",
            INIT_RAM_01 => X"DA51005ED2B2D65641D5ED47B9E700B4C02D987EAC05AA35452622C44020A840",
            INIT_RAM_02 => X"8208888A2A80EC6C6C6C5FFFA0464ECE00C6BF179558013AB820802041A020DB",
            INIT_RAM_03 => X"4F1DD430625D456997FE24653557F160F01FFE008C50A7610CEFC3008439C2A0",
            INIT_RAM_04 => X"8DB3DA83D40183A14B9640D09173C42045012C1B51100B8C664810CB08A588C4",
            INIT_RAM_05 => X"A2E903E7EB0DC011ADB3DF0D8D2376E69A630325200B96B0B628634B7BC40992",
            INIT_RAM_06 => X"6008011016DA6D04D848A45D000017972A89FF71E592564079FDE2C95590783F",
            INIT_RAM_07 => X"C05FEC0CCA1FE960AAC505410E4D0B678A965605BBA40A69CA97C8135AC04422",
            INIT_RAM_08 => X"83DD67FDF9F5B25C2D6B6ACA481827FAA71A0B0018CB4174288C92093DAC948A",
            INIT_RAM_09 => X"C5C2D9F623A928161080108EE344C931350A2845B5A988C69344528E89B021A1",
            INIT_RAM_0A => X"E4C49D81509C448984888062B24F49AC102231D0D12EA818BA199988D144B7AD",
            INIT_RAM_0B => X"012C0040C79DD38AC86EC13E5F18F0F12FA19049F88FD77C17241A85843AEC48",
            INIT_RAM_0C => X"EB10B8E6B47004A28FE8925F08F4375D0E4C1012A268F0222D88000A0DF5246C",
            INIT_RAM_0D => X"4AE58DAA300D44314D179A048E2CEBA48D622A8E1AA3C788D1E12C264187CE86",
            INIT_RAM_0E => X"56BB8380204A6762F1327228A521909845908849258C48F1D68C3511AFD652BC",
            INIT_RAM_0F => X"78D0777BFD10B2218171042FC0B500A0280C530771891E53E63786D55562A895",
            INIT_RAM_10 => X"2C3189369337D14258E5782ED18AAD135A5A1BA0F4ABF09D277428B846C66C18",
            INIT_RAM_11 => X"ACCC5F029EBB669179297916DB141336797F5AB94BEEECD7DC89E2C247C5AC56",
            INIT_RAM_12 => X"DE1281582A260159A225911041900E36BDE1BAA1D0F6395634543991B0A5BD8B",
            INIT_RAM_13 => X"B5495000012000608304141451E10A800ABAF507AAB3B62002CFAFA88B1BB82A",
            INIT_RAM_14 => X"80160108059B749002B490096003E6227003305A02B00DA1A0208B11860D5D5D",
            INIT_RAM_15 => X"AEEF98E268430B4D4220201234740EC621D0F4A28012600805829131830563A9",
            INIT_RAM_16 => X"0000000030050600002586259758B469047130012D60510415EAAFCEACA45408",
            INIT_RAM_17 => X"000000000000A2660788243E10B82800440000E00C4628100031913113000000",
            INIT_RAM_18 => X"CCC0F1D2449028A880A82AA2FEBC021C2FEAAFE64AAFEAFDA8197168045088B8",
            INIT_RAM_19 => X"80C3C8B6419ECC5893AD34912CCD27CB169EA866188810C01602220597202444",
            INIT_RAM_1A => X"44DB6DB7A146CC1A7288FCFD390D36EFC1211FFCE98398425B307888408ABC11",
            INIT_RAM_1B => X"997F7EFDFDCB310E411B1C01B4846DB6DB63B32C996E80E8910A42D386496A41",
            INIT_RAM_1C => X"2F112510C9555A484412393BB15B7C401D134F89B30CCC3D458CB237E5558CEB",
            INIT_RAM_1D => X"2E9323ED350D3168DB4EB5E05190FF573E0200F57D181CF8AD5A7A92A1811244",
            INIT_RAM_1E => X"6F34479DA3169899E821E9344786FFE2912FA9FACB21C62F6CD511F3D18DB249",
            INIT_RAM_1F => X"D929BE5019222E6C3FCFE7480D53DF6770F1328816F3C7290042AB20D992C84B",
            INIT_RAM_20 => X"5C8210EAEAE1F90284984B5857708B662A262EB6EC758467359164DB0811298A",
            INIT_RAM_21 => X"02EE2C37601024A058B2486BA1024777836E0E28152BD5FC192FDEB8F885FE30",
            INIT_RAM_22 => X"D42801000023773B6040D951AB0207400EE782A24890FA4818BAD86EE1C7578E",
            INIT_RAM_23 => X"8846B42AF82580100328C0417B875C1FC2DDBA37BEABEDB2850B9E9C40222D44",
            INIT_RAM_24 => X"8A600C8222278E4214844E31800062100F4B89B4080F12B312240669A70D1F90",
            INIT_RAM_25 => X"2D8968AD5A1094BC6110BEB60D50A0259B58621085B80480132C23EC294E4394",
            INIT_RAM_26 => X"3C28D04820A795BAB1983001B35E78E399B39AE0C7EC70E60032DFB9CCF95011",
            INIT_RAM_27 => X"10A1BC810864A8C020A2870F2A9D40EAAD1898A88EB885B66B9E8A71896CF630",
            INIT_RAM_28 => X"56640D839D332326E0830826B7AACDF519A4A9055920408820A66800408A7483",
            INIT_RAM_29 => X"20C60E789174010000622AB91448015B0C00696849C1515600C204586C046B30",
            INIT_RAM_2A => X"82DD6D8820942A05D30440E809F414100010DC84D75EBD2802288724B5013913",
            INIT_RAM_2B => X"F54C59C40966C393AA54BD63F03434E2307A51022074036D85233AD02A7E988B",
            INIT_RAM_2C => X"098528E097E27B124D10AB64DB76D48007276DEC0116D69F87406868413F6B28",
            INIT_RAM_2D => X"11E83C393E604EE855484C778B176497DE5012DB99941A985A6336450A929630",
            INIT_RAM_2E => X"28A4CBB0735B8D4B65D0468D216620FBAF7B0D4144021F842E00102420C04620",
            INIT_RAM_2F => X"B877683FC308E94E89E0AC24313A783130A4402D1102852A886D827731E59409",
            INIT_RAM_30 => X"99058D53FAF5799DDBAC36CD01F578C9146317AAB59E917FADA54727A93FDC13",
            INIT_RAM_31 => X"F0954D12089D460E96C834BBDCF7B9CE67318EE26C6D084AB131A9F814591215",
            INIT_RAM_32 => X"58FA75542203B310A2C6E6AB30915214BD00C53C40328A5E20BB3EEE80197D53",
            INIT_RAM_33 => X"212B9687395462D5522105E1B20509E88FE28002A3698983F7B3C4A875484416",
            INIT_RAM_34 => X"CEE9BD366E4D67B27593EACED57F9EC2C1D824B4F3002110B20E6CF4AA8705BD",
            INIT_RAM_35 => X"C2394768B66DE6C7C5DAFEF1186FE7BEF9BE6CF33461B0BDE3717A491202BCB3",
            INIT_RAM_36 => X"E4DB6DB42C8231F8F67B3D6CE971DE79325F9A64AB1D2FEDB698F5BEEE99370E",
            INIT_RAM_37 => X"8ADFA22245AF9126891E2245588A17DDD844A800963008732CCB25E69B19138E",
            INIT_RAM_38 => X"0721380F3C479CA1BA006B28665658E8E9E67E0010B00024B7372098EADDB8DF",
            INIT_RAM_39 => X"5374CA9AAA94C88B98008183373F959DF936C7632151B67642749AB949747BD4",
            INIT_RAM_3A => X"CC55A7674A56AE1767DDB349FF33EC68B1601E2CCFD73F88A9C3F251D3622E99",
            INIT_RAM_3B => X"DB7E95E739DED5F6E37BCEF381254E2FCD301103E960B26891A4480AD168F97D",
            INIT_RAM_3C => X"B8CAC5A2BEEDDC1DCE5EEDB9E07F76CEFFFDDC6FDFA8AB07F7FEEEF7EF775555",
            INIT_RAM_3D => X"283026E51A68842408A0087186243C800A829601D5842C0700D1401240CC6516",
            INIT_RAM_3E => X"47C93FA0638A7D47D23E2F1D80760060EE89142D20687BA55FA4A6595C011000",
            INIT_RAM_3F => X"FFFF000000000000000FFA33964F89E7BE76BA9FDB5DA9F6ACFBBE3FB9DF49F1"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"C1DE24BCE20FD7D600007FBA5F68BFFFD3803E5EEA7F940636A4A40484841C57",
            INIT_RAM_01 => X"7071407050EA52F7B9B9BB0EDF1F313C82ADD8DCAFFA0CA1952943A000103838",
            INIT_RAM_02 => X"2A0282820888EC6C6C6C6DF85E121612001EE2099948001A1851317141705051",
            INIT_RAM_03 => X"5D7BC7B9949D929516DAA5541016D800FFE000002429EF232BAEC000ED3FCAA0",
            INIT_RAM_04 => X"7977A4B0259DEE2843CBD6A02273606957A1B780153A02593ADD3EEDDEF7C0E4",
            INIT_RAM_05 => X"C5F22FEF939BA4412923C5812AABE74001602BB67A9FDDFCFF2F7953FFCCA1F9",
            INIT_RAM_06 => X"0008031020410CEAC0DDEEF14554545FA840BF7BF1E2F6CAFBF5C8F19DB3FF3F",
            INIT_RAM_07 => X"208925C8080927F8CCA1004B9FDDD964CFF38EE0CC912B08F8C48ABA5EC00120",
            INIT_RAM_08 => X"F7D53248BCF592D1AF7BE3004501F248BADCFFF760BB08442000C340192F30CE",
            INIT_RAM_09 => X"70745ED7B53C32ABBFF0FFFAF951217D1C232E047DE9E08693F0C08F1F75BFA7",
            INIT_RAM_0A => X"82109B494A0570E1A48F6003BD4BED2F803482FC048B0E4A9ECDDDD2FD123470",
            INIT_RAM_0B => X"808C2AC460C440BF8FD5CDFD0DBA7DFC2B83D8E53EA755DF1BA418C72048270A",
            INIT_RAM_0C => X"E2969DC57D1C00B08F7AF3175D333A564FDF455638B278600580289688E747B4",
            INIT_RAM_0D => X"78D581E384097199080A0A00DA47B69316A1A6DA97B424ED0939AEA57BEF4AEE",
            INIT_RAM_0E => X"4CA4C2529F5F25941B264BAEAD6B55A5C7C6BA49AD0F4D513E9F714145F15E30",
            INIT_RAM_0F => X"ACE8240E5F5598EAB85473AA80B02424A82053113183CE6C439EC4B33E66F905",
            INIT_RAM_10 => X"3EAB9B60FFF1FDDABAD3201055EFEC5E7EF63FD0C62B1000AFD67D7DFFD554DB",
            INIT_RAM_11 => X"940D4E82E68940B07A200A0A3BB2088508C7099AC320AA4C850020474B0052FC",
            INIT_RAM_12 => X"11528856EFAE34C10AA4D4E1C3F41A32B7837B308191911A242020E2943A4F7C",
            INIT_RAM_13 => X"3C08456416440000C201062818A1888008BDB9021BDDDABF2E0808BEABCCCAA6",
            INIT_RAM_14 => X"F50D018034AA75444624B50A4803FBE76800981203A009E3240005FEC4035C51",
            INIT_RAM_15 => X"BAABDAC087280BCB082A82056314002209C070080242010287E795DEBD67BC6C",
            INIT_RAM_16 => X"00000000000000000000000000000000000000000000AEAE45FFFAB5041F940F",
            INIT_RAM_17 => X"00000000000000000000001C0F00100000000000002000000000000000000000",
            INIT_RAM_18 => X"66400000600000C8080AAAA07CE6BDFB3AAAAFDDFC0E841347A3315588210040",
            INIT_RAM_19 => X"408B6F9ADBFFFEFFFEA1D7FE007A1BDFE1D7387D12510BFD1E4000903F200104",
            INIT_RAM_1A => X"FF5864EC7FFBF13DAC5FD60DE01FF8AC9039F337BD2442D7FFF82E7860AE9BBE",
            INIT_RAM_1B => X"880378F1F5587FEF4B5AB7E1FFFF6FF8BFFFEB4BFFFAE12FEFDE7D030810BFFD",
            INIT_RAM_1C => X"AC052868C53F52DF8A3E4AAE17C903F030F703AB0C39DE766C7AFCB39F71EAEF",
            INIT_RAM_1D => X"6BBFD5F01F0FFBFEFFFE95A043FEFA556F91C368025A59DF55E3FFEA2364425C",
            INIT_RAM_1E => X"8D7FA1F510E96F01BF900502FA1744F90AC2D607057FA30A61FF172045001000",
            INIT_RAM_1F => X"9140B47FBBFF8460B5AB4C2915895EF889C0D43A72BA75D7F887B6C91CFAC85C",
            INIT_RAM_20 => X"593ABDAEA2AFDF32FC9CFBDECD63DEFAC3164ADB480031A57C9FF8E03FAE1053",
            INIT_RAM_21 => X"91BF987A2BB6697872F3DDFD39F72BC6816B0B9CB57961D9CE5CF7AEEA2EEC62",
            INIT_RAM_22 => X"F1D6BE1111AFDDE15836B6A8F60010775C0E819ED524C9BED38780F425A3E6FD",
            INIT_RAM_23 => X"F3F07B49492D50112ABDCB497FF99D0A327117B9432A85FC40D83DF1FA0AD3F4",
            INIT_RAM_24 => X"A07D22ABCAED2CE3BCAF624A20A3BFD05188F5F4F80EC22ED03903C9E6CFDF89",
            INIT_RAM_25 => X"EFAB288C5F1FF580295D87175245CF03555F1CFEACB015FC57E9684F214E631C",
            INIT_RAM_26 => X"F7E03EF6FEEE2F6CFFE27807C9B3C33232CDFDBD76BD9632006626B14909F48B",
            INIT_RAM_27 => X"87EADBFA39F33EF17693E659D59FFB533E94FAF88BF74F8D1147F5F7BFDF7BFD",
            INIT_RAM_28 => X"CFFF9BD345EAA6FEC8A01350FA0EFEC9EBEDBAAFF7138BBB4C90FF6037BC7E79",
            INIT_RAM_29 => X"95ED1503BD40EBE764DCC443F59F6FE290F570E7B6A2BB2DC1BA8F3E8317D7FC",
            INIT_RAM_2A => X"26964182B2B3F681436E93C06C0922603BB05FB86EA53A11F69246C88A233633",
            INIT_RAM_2B => X"A38FE0FB6618A00FF07BF2C900787053EA76DF2EBD835041D3F02AA2615B1EB9",
            INIT_RAM_2C => X"9B1E791D13BCE9F2C249A965DB76D69AAF21FD163577FECFAC830990D577C232",
            INIT_RAM_2D => X"098757837ADE4C2A30E05DAE56A036D223FC8FE37F7D0131FB6EEFDFEF9F3D0A",
            INIT_RAM_2E => X"ACE6FAB4773B0FD36984CF2F6BEE2EFFC7781B937DFABF2867EC1E2CF8CD9D35",
            INIT_RAM_2F => X"BB7F5AFFFBBDE98F138D2E7DBA7CF13A706C8A89001489134C59877F63E9C72D",
            INIT_RAM_30 => X"F51FCF7A5DFDFFFFFF9CBFDD45FA7B9D346337593D9BA5372FBDC727AABFDF33",
            INIT_RAM_31 => X"F0FF5DB37E9DF77F86CB3CF1CC639CC66739CC726C0D2CCAF5398FF93D7F561F",
            INIT_RAM_32 => X"5CFB17AE07ADFB9DEBF5D4FF70F5FE87FDD2E1FDF4BBC3CEF8EBBFCFCC9EF6DF",
            INIT_RAM_33 => X"35E586D155EF72B5426BD7B9FDAFDD09DF55B82B9DE3A3AB7E7FF7BD37AC4F5D",
            INIT_RAM_34 => X"8B690D264FC9553FB7874ACFFF5FDFE3CDF9BCF676070550F21F6CD7F2558B61",
            INIT_RAM_35 => X"C339D76AFE7F7F97E9DAA587BCDF0508AD334C9A3445E2BE8BC57AF9125AE922",
            INIT_RAM_36 => X"BFF864BA6FF9EBD8FC5A2DE4687B31CDD3FDDAECCBD3AA79F5D5F1EEB6D9BB6D",
            INIT_RAM_37 => X"ACD26AEBD5873503AB58EBD579AA05D49808098EE7F46EF64F9BF77FDBDA3E5C",
            INIT_RAM_38 => X"8FA1502FB857DDC9BB54C233E414196968654600000400002B3834DDBCDA38D9",
            INIT_RAM_39 => X"525EBA9110602AAB980183816B36D39DDB36ACD32E5BB64E5B2686FC587D2BA4",
            INIT_RAM_3A => X"F6468F667A96870736E6B31BDAAB684952A01B3CEBEFB9CD8B6BBB3BD7136BD7",
            INIT_RAM_3B => X"DB75ADE739DEB5B6E77BCE739DE74E7EED76B3574B47FB7E9DA746EEFDFED57F",
            INIT_RAM_3C => X"010107EBD7AFE3E3EE5EEDB85777B6EF67FCDAB7BFD0D0AFFFFDEEEFEFB6E26D",
            INIT_RAM_3D => X"0200000080040A004400440048008010012000A00040028009000100090080A0",
            INIT_RAM_3E => X"5F5B7BB67BDEED5F52772D42D90B677B88A33517EB50222D57BFEE0204040210",
            INIT_RAM_3F => X"FFFF000000000000000F6AE7DEDB8B76ACB4F3BBDB5DABB38DDB327B49DB8BD8"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"17133C5624CAB161000CEE844AB02046428CAC32B7CCA2CBA1A5A50D0D0D1D71",
            INIT_RAM_01 => X"8F8E018FAF9909C203D688627906C86195716CFE5E0D796D2C04805F7FEFA8E4",
            INIT_RAM_02 => X"00AA802A0282800000007DFFFEDEDFD200D6D201080000040220C000008021AE",
            INIT_RAM_03 => X"0639DCE7F6DA35FFCE683044FCCA41F3000000019FA88CE67E7A7C0198792AA0",
            INIT_RAM_04 => X"49F381990CCF222B5F00591389ED02C046707409A1E706037633D39D398CB599",
            INIT_RAM_05 => X"31CCC3024E79C758E59B24E58422311B2C97BE5EE548349A90BCC00E4E110D84",
            INIT_RAM_06 => X"E4086132596486332CE2510320C31C10888BA4C08F1A0F7C20971F8D63DE21E6",
            INIT_RAM_07 => X"40ADB658E26DB566AA922A334A75077698B7E36EAAC98425C3DEE660294B1886",
            INIT_RAM_08 => X"98C4AB688F7037CEE529062F28FFAB6CDB4C433558DD25C064028A2CF90C662A",
            INIT_RAM_09 => X"41491846616425567397F39363732771BCB0380A3286865A4BA759A64912611A",
            INIT_RAM_0A => X"793209037B0DC38EB2DF7206136320BCDBE040D31D32396B3BEAAAA1D374DCE5",
            INIT_RAM_0B => X"7794B9DE40E45CF84520470C7C1B10C19D9080D1B9B71F1C21B24BE96C2B0667",
            INIT_RAM_0C => X"C61DB8E4127192525B23987BB83A2064B65C61E6E1B45BA6E6BD9BD0BCBC2280",
            INIT_RAM_0D => X"CDE2128E2009C733268409378A44A29AB4718F8B12E0049801241444C3852E82",
            INIT_RAM_0E => X"FCD0CB998F7E25C075EBD8B1B5AD36984DCEAB66BCB578519264938904423301",
            INIT_RAM_0F => X"F1841498E0DE39824588C8934033B336EDB8CB21079F1AC32A3DF7773FAE7FDC",
            INIT_RAM_10 => X"EC10EDBAD339904BB14B7208DB2299004A32D98B0E903029B26D6060664CCE08",
            INIT_RAM_11 => X"7704EE480FD9D4B8DE4C0579B309EC4D8EC76D9CC599316CEF2C250839180B35",
            INIT_RAM_12 => X"24CB1C339B9CF1E41B369EF82D81FD65301905768293F73A6DA0E46EB2E22C3A",
            INIT_RAM_13 => X"25E420E014001800C0850E3031B141000136310E66F15A26DF22816E462AA89F",
            INIT_RAM_14 => X"D08C653DF2ECD74DDFDC53670403E666E4F0513ECA95658C02F39732CF793F62",
            INIT_RAM_15 => X"DBC9BAB41507030B6599D9531124290641996641D9394890CD86070AD5B4A4EE",
            INIT_RAM_16 => X"00000000381FFF00003FFFFFFFFFFFFFFFFFFC01FFFF041011FFFFC050555009",
            INIT_RAM_17 => X"000000000007FFFFFF8E3FE3F0FFEF807C0000E07CDFFFFF003FFFFF1F800000",
            INIT_RAM_18 => X"EEBFFFFF9FFFFE0A820A28A3FD14414D2AAAAFD4500000401100740077DEFFBF",
            INIT_RAM_19 => X"0064D4F181AEDC1DDA7386D0004CC1830345506C5F73197AD41F3E67DF90B7B2",
            INIT_RAM_1A => X"7C35D784654FD77A773DB9BBB76D33925871AF6630B3390F0D30610C5312FA7A",
            INIT_RAM_1B => X"A2AD1B17466DB93824277B3324C4DDB1D36F210C99738F56FD23CF2F65C8AE02",
            INIT_RAM_1C => X"1F1C90F3C5BCDBB99B3A26745CED804D1041BE1884280C07FF6672391CF13E67",
            INIT_RAM_1D => X"F87348E2459DB079D26DCA809F930B45B6E849A5C7212449A6443FC4D3BFD932",
            INIT_RAM_1E => X"161491D34964B92E99D807DBCB8676CE6EC58663C1F59277F6F112BF33FE0800",
            INIT_RAM_1F => X"C69258900F3761B6341355BA47272DEBE45B1EEDDC71C32B092E7F7349957814",
            INIT_RAM_20 => X"226442C9828349D93329652B7418B8E25A4F9852711B933DB27BB3659D66C820",
            INIT_RAM_21 => X"29CE81919E6BB42010A65663E78A910B1ED8087848211B4F34891A61E110A7B9",
            INIT_RAM_22 => X"C7ED4037739677A4E20CFB44204FEF9C879B02EB49BAE75B00F3F32392110B0F",
            INIT_RAM_23 => X"8713F96F4893A3B6D60B74F5888F7EB604CDFADB8C2267B164265ED3C8D9AF72",
            INIT_RAM_24 => X"E5BA59EF67BC9D5ED3B6D964966FA64B38669997EC6819E65BE6806DB76C1CE1",
            INIT_RAM_25 => X"B69D6F3118F2D660B46808BBADFABE844D1C99F2D27E3799DF1A97F4E73FDF77",
            INIT_RAM_26 => X"3BF7F3C0679FEDBA37AF709F3457E10C0047BBC6DB66D27E00AA546C26271875",
            INIT_RAM_27 => X"4D8EDD8D90EEE5D4C02E5A27ACE549EA8CE7C9AA0A38759485224A10813D3673",
            INIT_RAM_28 => X"5CCC8D2A27B12B6642946D89E7384967AD802B1D78EF766C3649A9C8879B7227",
            INIT_RAM_29 => X"6A9E4EBEF1C135CE9BEBBB233739B76F6C5ABFFFFFDD445E83D2B5FB84C44F73",
            INIT_RAM_2A => X"4BB0F3FDFBFBAB3E70AD28D63E365DDE35CC47674746FC84E9659F1654CD59D6",
            INIT_RAM_2B => X"CD3DD0DA90FE1E692C7095E50033185E61A37198779FACF2AF0CE1CC98C86EE7",
            INIT_RAM_2C => X"6704A99A6ECE312B34B2EC9324C93D856C9D27310B9AF278FCE825696A9ADAC5",
            INIT_RAM_2D => X"C2A69FE51C292DAFCF690C6213CF692FC65000EF191608501872306542C256F1",
            INIT_RAM_2E => X"99BD4C5BCFE6796DFFA16248B726264E0460C02DC61E4716161733B3B68776F2",
            INIT_RAM_2F => X"61C4FC310E699838CE08F9ACE1E3C0E1E2B795450023A74F88C186C46887188B",
            INIT_RAM_30 => X"367734C586F12919C969E6430499CD7E498C4B00373ACA6CF8663CB67531319E",
            INIT_RAM_31 => X"F09104E2E9F2048A59F9E3A5295A52B5F4A56B4B58D6A679A1A6B8F872C99071",
            INIT_RAM_32 => X"638D8C630E518273964CE0890893125C3D07973F41E62E3FA0844A3B267275F1",
            INIT_RAM_33 => X"55245B68131C4ECAAD7F2C25CBFBB303476F99767726E6E3B1F3CC938C761CB0",
            INIT_RAM_34 => X"2EB2464C9E9366725C85BB349188481E5CCB8F93CD81F11F92C4B6EE800487A0",
            INIT_RAM_35 => X"12E371B5D9742632672DC0810A070C49D67598AC91D4EA3289C467C6C5CFE20B",
            INIT_RAM_36 => X"B4D5D763398461E2712C972137CF6797255E6D19D670D2431A7059339B792DCD",
            INIT_RAM_37 => X"CD6AB8B972D31C2AE1CAB972C8E2FE7B8267E6414C90941DF97E5C266D345A04",
            INIT_RAM_38 => X"9B2B9364E3723016DCAA9AC4764663B3B3B67B7F7CFBF9FC60D80C41DD685368",
            INIT_RAM_39 => X"AB6BD55C0460088E5AAE8EE1349B3E43450C1DB087FC9921CD1A632843CE8289",
            INIT_RAM_3A => X"3BBB7C91AF88AEDADDA6CB19EA23AD72A54DECF21D1E77C41182CCB0ADD10D7A",
            INIT_RAM_3B => X"3B8B93E8B9C07662E0F8108C1C1DEBEF368D45A9B99E92EB76DDB3D947234323",
            INIT_RAM_3C => X"FEFEFB278C9DFFFFF7E31DC7B788231FE7FFFEFB7FAFFBAFF7FFEE3F8836E76E",
            INIT_RAM_3D => X"FDFFFFFF7FFBF5FFBBFFBBFFB7FF7FEFFEDFFF5FFFBFFD7FF6FFFEFFF6FF7F5F",
            INIT_RAM_3E => X"C12F2853CF3627C13D1194604DC133C998A19D826C89D5A7E364827DFBFBFDEF",
            INIT_RAM_3F => X"FFFF0000000000000039261E7272891A61DBED8924F27899DC4C632906E9BC42"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"328B18492E490203000DA28440801002C24CA434B280B2CB8381810909091923",
            INIT_RAM_01 => X"00000000014909A0065259257906DAC195417AC95E0A29672C4D8000000021AC",
            INIT_RAM_02 => X"AAAA8000AA807FFFFFFFFFFFFFDEDFDE00DFFFDEDFDE00DFFF860E8600078600",
            INIT_RAM_03 => X"0A3088C7F25395FFC90420447DCD2800000000019BA808E6FC3534010C40000A",
            INIT_RAM_04 => X"49E12089044A227BDA005B13AB460060CEF0D00943EF06084477811410529F13",
            INIT_RAM_05 => X"7107E20404784758CC9A64CC8E2251092D90BC7A42456C08A8B588040C3B870D",
            INIT_RAM_06 => X"810001325B2D863364EAD56371860C11808B80891E1A480E41123F0D720240C0",
            INIT_RAM_07 => X"2880029802524A051132AA6E1C32082811B4048D11318C6C8B9EEEE1719B1A84",
            INIT_RAM_08 => X"1B22000187682DA19084066769C380011840483100102488E4668A6CED403353",
            INIT_RAM_09 => X"010C0000601404006017E31981768EC19D94002B230E04DCD9E31B653021053A",
            INIT_RAM_0A => X"833600037981860F36DF1235036629B8C9E060A20C18313195F33331A23068C5",
            INIT_RAM_0B => X"13B99BDEEA508A78452087207899C1E5BF399180E1929A307192C9EA6C63C56F",
            INIT_RAM_0C => X"EC0DA800212096D25C01107B18022170183035FC434AE94EEF1DBBD394DC2280",
            INIT_RAM_0D => X"8002170C28088732648601338040A01B34018D848060A01828063440A6062504",
            INIT_RAM_0E => X"FCF1DB9BAF3E26B0F5EBDAB8B5AD16985D58BB2E99B9780000E0A61804032008",
            INIT_RAM_0F => X"900415B421CE3B826DCDD8B2682397166CB9C922073E0C40281D6B777FA67FDD",
            INIT_RAM_10 => X"E810EDBAD32E800B918956189A201900C932D91B1E811821B029404066444810",
            INIT_RAM_11 => X"F3E4E6C52FD9EAA4EE440F7B151B27988672B49E663B9B2727242548790A1B35",
            INIT_RAM_12 => X"65DB1C63999C71EC59961EF8288154645039073202A1F33A6480A866B6C0383E",
            INIT_RAM_13 => X"20EC69E8040C0070C18102380882E98809B9790CE66124068F628166CE1110BF",
            INIT_RAM_14 => X"500A251DF6EE634DCFDCC72F0E30D8D01050C33E4A9727064673B6224F396B37",
            INIT_RAM_15 => X"35143425350C861B2CBBCB9D8CB04B4E53C92251CB7B519440154692D5AA94C4",
            INIT_RAM_16 => X"2110921148211104104108889042052244844412484950101400001500554186",
            INIT_RAM_17 => X"22222224924892492492493D3F12209084204920854484211042221120822222",
            INIT_RAM_18 => X"888000000000002A880282820040411015555005400104545111441710422489",
            INIT_RAM_19 => X"006434C988B25425491692480024C284830CD02C4F331988700000000E00B510",
            INIT_RAM_1A => X"0A2CB7A0540D536A7735EB96B769219258D0AF6294B1391D14B0530C37347AEA",
            INIT_RAM_1B => X"22251192A328A8A5242568969442B4934921600448134F5010282F6764C88663",
            INIT_RAM_1C => X"189DB1F384BCDBF5992A2650CDB680201052350884240C0FBD6A22619DA1A222",
            INIT_RAM_1D => X"F169592245B490B5C92BDA40CE8B0944B4C041A7C7232485030E254E5AB5CB72",
            INIT_RAM_1E => X"1A22B3535904B526D5C802C9A982292E26C180EBC0D5327356B002D3338E8800",
            INIT_RAM_1F => X"A392C8A0169561D262395490CC2CB5AB848F3EECDC51A282092E7D733B978014",
            INIT_RAM_20 => X"32EE46F44743A0CB332967797288B4804A45B452F90B971CA26A91AC95664860",
            INIT_RAM_21 => X"295A81A3BEE9B410108D5212C698B29D00B504F8409089A724891D115010D3D9",
            INIT_RAM_22 => X"A644003773B732ACA20DEA0C8240000DABBD02E94898E71900937347B2329D0B",
            INIT_RAM_23 => X"0F43A96709B2A234400BE0E1850D6A384EA5E8EA9B226293242E525228F98636",
            INIT_RAM_24 => X"ECDA59E567BA9B5E5396C92CB6EF845B796E195784249BC45BC4022D142A1265",
            INIT_RAM_25 => X"590D67B514600241FE288BAD05F038045D1499E2D22C3719CD12939CEF39DEF7",
            INIT_RAM_26 => X"23F3AB80411E689A10A7508F3057A10E1086AB568D52821400AA44682564B876",
            INIT_RAM_27 => X"DA45254D90AED754E0214267840409228464CB82010820818F65402108B51553",
            INIT_RAM_28 => X"5AAA84AB67912156C2946C9955340522A5A48A1829ED22E432D9C5D8275B6AA6",
            INIT_RAM_29 => X"605A0A0EE1C100DE1BABB9662771B0250010DFF9F9441C5A8152B0EB82440D51",
            INIT_RAM_2A => X"CB68B6DDD9620335928D28D236B6DD8801DC0B3741445C84E965B912404D65D5",
            INIT_RAM_2B => X"4534505AB0781E6B8C31A0A70037285161D32898D79F85B3068CD14498A47666",
            INIT_RAM_2C => X"2304A100375E502B34B2C6B36D9B6012698D4730059A7420FCC00441522ACA65",
            INIT_RAM_2D => X"43002FED142B78B3CE650C4411C74DBA564010A2191004701052364442C25049",
            INIT_RAM_2E => X"19BA004287E6516C9FA364DDB740040C0040412CA2064B160C3303B3B28376F2",
            INIT_RAM_2F => X"40887620047B1071C50071C8408140C0A080D5610031224488C1028859021C8B",
            INIT_RAM_30 => X"B6729ADDC6EAA485D569468600188D36CB18CF0A326A40E650C028B67F20238C",
            INIT_RAM_31 => X"A00A88B163204D894B0943AD6B4AD2B5B5A5294B4C88623503EF90D02921126A",
            INIT_RAM_32 => X"F70F4263042146E1490C285A1802A0482805122981456414C046C933222220E1",
            INIT_RAM_33 => X"74044BD41098DC4AA95A12875BEEB703C92D182976A6E6E6A8E10A5382760848",
            INIT_RAM_34 => X"26B646C992B232485D159B324A00003E98530BA10C85F11BA2C8B7AA544D86A0",
            INIT_RAM_35 => X"326721B149D202606231518112448C44565598ACD3C0E022A1D047C2448FE309",
            INIT_RAM_36 => X"12CCB7C3114C41A65164B343128E2592245A6C3BFC70F9229870889199796CDD",
            INIT_RAM_37 => X"C58A90912351080A40889122D042FA6B866006D318A1B04CF13C4A023170EA08",
            INIT_RAM_38 => X"B92A5340C1606096E0AA8A6452C2F696969329000000000060E80A2155886388",
            INIT_RAM_39 => X"A93955491060088CD2AB0EE015897EC74C1C5CF183FD1B23450A2130068EA3A1",
            INIT_RAM_3A => X"3BA955B0A588AE5ADDE6DF19AA22A536AD5FE5F6353CD2A200A24DA52C88872A",
            INIT_RAM_3B => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFDE9ED361D4DA9999AA2E932CC9155A351A706",
            INIT_RAM_3C => X"10001B858E1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_3D => X"0004008002010040000800100100080020002001000800040020200100200004",
            INIT_RAM_3E => X"422D10F28B7646423F20B870C5C3128899E089862D89C4E28062040000004002",
            INIT_RAM_3F => X"FFFF0000000000000030020A7417001C01C9659124B25919CC8C43110F70AC82"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

end Behavioral; --VZROM
