//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Thu Dec 14 10:24:48 2023

module VZROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [13:0] ad;

wire [30:0] prom_inst_0_dout_w;
wire [30:0] prom_inst_1_dout_w;
wire [30:0] prom_inst_2_dout_w;
wire [30:0] prom_inst_3_dout_w;
wire [30:0] prom_inst_4_dout_w;
wire [30:0] prom_inst_5_dout_w;
wire [30:0] prom_inst_6_dout_w;
wire [30:0] prom_inst_7_dout_w;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h9E2AC9857A68EAD3001FD1BD57A9D4A75B240075E080974B999B990B092B1923;
defparam prom_inst_0.INIT_RAM_01 = 256'h179AC0C6955DA9AB53165DA56082DD5F3FC55F63FFFF0560AE9E8C1EF4CD50AF;
defparam prom_inst_0.INIT_RAM_02 = 256'h28A87FDD5F827FAAD50023BBACC88A5240D3B18D0EEA417AAD439592C1C294E1;
defparam prom_inst_0.INIT_RAM_03 = 256'hAA89185FF3443FFFDD655A00FEE50A9753F9B5A5BDD602E6FC9C7C0B0CD0202A;
defparam prom_inst_0.INIT_RAM_04 = 256'hC1126C1D60EAF112103A3B2B9802006483726829C0F724E1127B817A1118157B;
defparam prom_inst_0.INIT_RAM_05 = 256'h581EE01464F32798B495246696057138F5A2F5DD4701B99429FABDA5883B8E15;
defparam prom_inst_0.INIT_RAM_06 = 256'h870060B279A696232CD54A8724925956924782AC0A713C1E10029538CF0700C1;
defparam prom_inst_0.INIT_RAM_07 = 256'h98B7DDE8B07DF7BF675000B8A6954CDF790187DB6753D19E77FD776898AD2D84;
defparam prom_inst_0.INIT_RAM_08 = 256'hBA88DFBF6EE2878FD294969FF6F79DF7DE6E4DF7E19DA397F4936D2EE9B51E22;
defparam prom_inst_0.INIT_RAM_09 = 256'hF2FBFFFBEF563EABFADBFBD8B613F71C2AD91A49D994B705ECFFF890CBA2BD5B;
defparam prom_inst_0.INIT_RAM_0A = 256'hFD164D880F09EABD3E02224D1B613506E3CE835D7EEAFF9C61CC4C795DFBAF7F;
defparam prom_inst_0.INIT_RAM_0B = 256'hD78BBDDE977A5F73A7D08E772CCF1E4BF883A8310BDF198530FF7772F8971AFE;
defparam prom_inst_0.INIT_RAM_0C = 256'h3EE80B453BDFDB19D527F9F5539328956AC7E5D0F1BE2996E33DDBFA355D13D0;
defparam prom_inst_0.INIT_RAM_0D = 256'hFBF6799FD00AF266BB975BAFBC572F17C5E387BB974E37F38DFCC197D8F312B4;
defparam prom_inst_0.INIT_RAM_0E = 256'h7CE75A9B9BDC91F93A443BB80942206E9640F1B4BE0BB3CB7B6DAF7DFB61FEDB;
defparam prom_inst_0.INIT_RAM_0F = 256'h40BCA00582FF6DC0678CDDB11F1BDA3775BBEC2493BFB5FEAF6C7B795FEB3BD5;
defparam prom_inst_0.INIT_RAM_10 = 256'hEFDC425BE002BC8FAEFA96F70F67484CAF3B804E1E10256CD28A262600008F14;
defparam prom_inst_0.INIT_RAM_11 = 256'hF3376A4873E4FF0A7EBC933B2D59EECDCEAC6E4F339AA96A7B5CC69DFC1D27B4;
defparam prom_inst_0.INIT_RAM_12 = 256'h7BEB5CFF3DD975ECBFBF6E3D1A83818926314B174348F7BBE1D0FE2C9FFD141E;
defparam prom_inst_0.INIT_RAM_13 = 256'h03EEF6F50A502001C20210088086038003E7F50EEF7B4EB7AF7587777CEE6AFF;
defparam prom_inst_0.INIT_RAM_14 = 256'hF299BEBDFE62276EDFBDEB7F3623C00280D2DDFEFDE0B88DDAF7C9BB4FBAF7D9;
defparam prom_inst_0.INIT_RAM_15 = 256'h26AA686F9FA7A524E7DDFDE6CC2C79F3FCFDDF7FED3DFEFFCAE4662E3C78C677;
defparam prom_inst_0.INIT_RAM_16 = 256'h211092115827B504106A5DEAE29F59569B2688135B91155195BBBA8EF57DBE88;
defparam prom_inst_0.INIT_RAM_17 = 256'h22222224924F14F9C19269692B548E9098204960DD8B5DAD1058C64E24022222;
defparam prom_inst_0.INIT_RAM_18 = 256'h2247C2DCA4ECC89703C78A224F40BA5D2BEEEEE7D919BF1D4F2CFF9931843D0A;
defparam prom_inst_0.INIT_RAM_19 = 256'hC036D2FDE0705521007A28009201C20401C596298FB5399D2A5C6C224D00B612;
defparam prom_inst_0.INIT_RAM_1A = 256'hA877F3BDD6FD5FEB79B1EBCA3BC209AAB8F80FC894F2BD3C143803EC5F6436E3;
defparam prom_inst_0.INIT_RAM_1B = 256'hAEE8822485450EB1B4B563FE9F18F497090C69C50BD51C2D5AD50FCAB5E91CBC;
defparam prom_inst_0.INIT_RAM_1C = 256'h41BFB2FC1D8FC0F1FF23B7C1E6B8ABAA748AC8402E350A0BFD6C4E4ABD406D54;
defparam prom_inst_0.INIT_RAM_1D = 256'hFD6161222DF41471A98EA9406EA3A4AA01D4CD186FA7A6E158BB03137ABFFF7A;
defparam prom_inst_0.INIT_RAM_1E = 256'h8AA8C21B28D371E7D1FC5FF78CCA93AB38E4FDB74E44517C84379E5C78F3D926;
defparam prom_inst_0.INIT_RAM_1F = 256'h715F2B2F920421424048C1C7EABE108AD68F8FFDFD5582178B77FD774288A836;
defparam prom_inst_0.INIT_RAM_20 = 256'h9AE3420150428DDF3F94385618293144C1E2B114AFB8DBC20EE280B89176E9A1;
defparam prom_inst_0.INIT_RAM_21 = 256'h6912C4ECFE791E5031751A15461DC2B435D1007348C4B08FFBD00047115347ED;
defparam prom_inst_0.INIT_RAM_22 = 256'h2AD6BE3BFFF1BA3AA45C62B053D568FD17CC03BE2D0BFF3B847BB9D9FB428403;
defparam prom_inst_0.INIT_RAM_23 = 256'hDBA70BEE56BA27D56BDCEBA875FA93613B2A412A34D50293F4AF021A8D5BD7B8;
defparam prom_inst_0.INIT_RAM_24 = 256'h645ED86461D894240802A310976FB77BB9EED05BD670DDF76BF56302010200EB;
defparam prom_inst_0.INIT_RAM_25 = 256'hF386EFDE857B7743E6BB334356F57D4ED68E9DFA5E5F3DDBFD5BF9611A84B1A9;
defparam prom_inst_0.INIT_RAM_26 = 256'h0BF7E3EA779FFBF254BFD79FBE5FA9C0D556AB140453BE68000448EE77CC2B5C;
defparam prom_inst_0.INIT_RAM_27 = 256'hCF067106D9AF575F321957BBD566FF0C956EDDDE3C63FB9E9984158314B59456;
defparam prom_inst_0.INIT_RAM_28 = 256'h7AB890AF87C5EC469D52B5E854F56533F0109A3BEDF72AF5D7E8D1ECBB1CAA77;
defparam prom_inst_0.INIT_RAM_29 = 256'h3558E86BF898AACFED8FDB83A37DBAF45A353FF5F512AF98F115DB6B27CBAD54;
defparam prom_inst_0.INIT_RAM_2A = 256'h6D63FC7FDB675C7BA1BFAD5116366ECD0BDC83765C16FDDEFF759C774A1EEFED;
defparam prom_inst_0.INIT_RAM_2B = 256'h00B55C59BE3D5F4EC35663D20F2667596D41EAD9C78FD7F5563EC5E3FCA176FE;
defparam prom_inst_0.INIT_RAM_2C = 256'h76215115061E41B9B6BB4E9B24C92B5FF098337AFFF573747DDF1FD5FF23C035;
defparam prom_inst_0.INIT_RAM_2D = 256'hCD654FF8A17BA057FE78208585AE12457CAAC108020A892605000282C5342AFD;
defparam prom_inst_0.INIT_RAM_2E = 256'h1DBC042DAFE69767BF9E0D751E5C4C29021069AFABF72B5D17133B9FB7AFF0BA;
defparam prom_inst_0.INIT_RAM_2F = 256'h4088260024F215B16D4E53E049AB5349A3C1CFC480B376CCCBD40188090276C4;
defparam prom_inst_0.INIT_RAM_30 = 256'h377A6ACC0460263195045E724855AFFA49084043262A6E3B92421A4AEE0022CD;
defparam prom_inst_0.INIT_RAM_31 = 256'h0B032ABCFE6B6AC04FA149021215240B4A484290B7D0CA79FA15B184A38123EA;
defparam prom_inst_0.INIT_RAM_32 = 256'h1B05E8E3B47A15611C09B019C90620D802097601825C6C00C313547BB32E09E3;
defparam prom_inst_0.INIT_RAM_33 = 256'h5A4D497E2A38AD7FFF9A38820FEE7A4B47FD3CBC7E3FFFE4A31A0FDB28E768E0;
defparam prom_inst_0.INIT_RAM_34 = 256'hE493E278FA9EF7E1CCEC53702A80045E784F131BAC9352239F6BFD2D1068BEC9;
defparam prom_inst_0.INIT_RAM_35 = 256'h7AEE60D30A908721569109A0D340CDE703F0F287958080082110179B66CFEF3D;
defparam prom_inst_0.INIT_RAM_36 = 256'h68F7F359970FC10756BF1F3979AE79E2E480F4FDD5F7899269E4F847B7C01B84;
defparam prom_inst_0.INIT_RAM_37 = 256'h4A8AB0B0635F5802C580B0638CC7FA2B8E6556EBAB9FBB3DD775D8875172FECD;
defparam prom_inst_0.INIT_RAM_38 = 256'hF85BC642D0A168D421FF44341F467373737F7756194AB55C4FAE3C6E1E832A82;
defparam prom_inst_0.INIT_RAM_39 = 256'hF9697FC800189055AFAF5E424C807E63468DB8F087F9C9A90EACA3D019AF8DAF;
defparam prom_inst_0.INIT_RAM_3A = 256'hB1DD359ACB076EDE0C6EC9AD0E5027B7EFDDA3F3514324460034065DFD918F2F;
defparam prom_inst_0.INIT_RAM_3B = 256'hC08C2308B9DE71E2E080108C371DD7C07A7D77AC53FB9FF1B268D170AA548B94;
defparam prom_inst_0.INIT_RAM_3C = 256'h346628D6AB38F3E7CFE3104417FC771FFFFFFEBB7CF7F1AD77FDEE3F881CE739;
defparam prom_inst_0.INIT_RAM_3D = 256'h557E48B37DF232D3B2D5329E935F5347348F593A2D91D4A6F278B66AA26F3329;
defparam prom_inst_0.INIT_RAM_3E = 256'h022491E299FB47022DA088368CDA32BC444198751D95DD16817F94A49CFBA944;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFF0000000000000070801A25CD128057BDB691FE7F3D1AC68C4B906D516082;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h084738CFEF89F8CB0003043ADFD21DB81214E311121915C585838191B39301A7;
defparam prom_inst_1.INIT_RAM_01 = 256'h091900B66C77F23C83243194B9C5D4C39FDE77AFF20FEC5D892DA1D53688BBC9;
defparam prom_inst_1.INIT_RAM_02 = 256'h0A022A08A87FFFAAD50054A8AB449F9A00813B8BB04E006063C3031301B5E14F;
defparam prom_inst_1.INIT_RAM_03 = 256'h4F9091C00CB6680011E636C5821599E38952D9C6207E290082A4882C3412682A;
defparam prom_inst_1.INIT_RAM_04 = 256'hCDB9EEDD76C607394B9CFAC6037659A265014142991000ED54484700637B3F02;
defparam prom_inst_1.INIT_RAM_05 = 256'hF98BB6D5CC03C8511902D5AB5A37432713656C008F6799A1BE81894C14AA8933;
defparam prom_inst_1.INIT_RAM_06 = 256'hC4802210092DC022135DEEFB820809E0218A9B397E3A64B35964FF1DF92C5D9D;
defparam prom_inst_1.INIT_RAM_07 = 256'h70B7F8D172A6D7C2FFBC4033E41608BB831525DAFFDB3DFA8650822832929424;
defparam prom_inst_1.INIT_RAM_08 = 256'h0B19CDFFC186A01F8E738360002C0DFE68A68E0080360841180524430108F14C;
defparam prom_inst_1.INIT_RAM_09 = 256'h2927EFFD07DC43FC2C34AD3809FFE16BB87B5011ED3C1BF4BD50D1ACD0A7C7F8;
defparam prom_inst_1.INIT_RAM_0A = 256'hFB5E9644E9531F0965EA4801E5D25A719E27F729C11D2431B21DD54E28046041;
defparam prom_inst_1.INIT_RAM_0B = 256'h0073A83553BA071145A6016821802A1D21719EF3B0697458C4BCB85399963B48;
defparam prom_inst_1.INIT_RAM_0C = 256'hE82CA1E8AF4031D69C580B42E9DD4C38ED582F440F97E8CD9D33061891C062C4;
defparam prom_inst_1.INIT_RAM_0D = 256'h24082769000023100B33F4401E8A07A1B0B0481DA387F841FE11F4987B025704;
defparam prom_inst_1.INIT_RAM_0E = 256'h05B5FE96024099796B22DC68F6FD1BDCF9F0BC9C27EF01B825E0248626370955;
defparam prom_inst_1.INIT_RAM_0F = 256'hCB1815B79610D8F22E47105F7E7E002C0262158018707C8020D9900048109032;
defparam prom_inst_1.INIT_RAM_10 = 256'hA6DC8B322634E9A442F4699CD42F7B6A77E839E061F13C8D24126E6EC4444864;
defparam prom_inst_1.INIT_RAM_11 = 256'hD0B1111C6C0C36BB2123268345C4D3E21136C8C2FAB4EC934C83736383641C41;
defparam prom_inst_1.INIT_RAM_12 = 256'h9D06400084A0061386A501E742F0934D72C052A929078C81964A457A6094E9F4;
defparam prom_inst_1.INIT_RAM_13 = 256'h201210284A483020038A140031A54E800EFE6A0321056CCF788C4F1238F7FB20;
defparam prom_inst_1.INIT_RAM_14 = 256'h5780BA233405EC31100230484003F96F88E002C0341D852B00802C4D208158B7;
defparam prom_inst_1.INIT_RAM_15 = 256'hAA445B7124880256040810B8CAF41B49924471162040D0655A0C9CC0DC9199FF;
defparam prom_inst_1.INIT_RAM_16 = 256'h00000000080B2B000015D9A29C6ED6B604080401497AEBE7FB050450403B9D0E;
defparam prom_inst_1.INIT_RAM_17 = 256'h0000000000044978CE8432E75D170300280000C06892ACB100108EA60A000000;
defparam prom_inst_1.INIT_RAM_18 = 256'hAACC7ED8263EFF1FCBF00D67423CEC450514142FBEF873E0F99B50050148B8AC;
defparam prom_inst_1.INIT_RAM_19 = 256'h001BA01B88A173076DEE416D25B64EC0C4476891BA005DC79C13024797002566;
defparam prom_inst_1.INIT_RAM_1A = 256'hF9E2083FDFF1202508936634C80F3E73F150C6010E668671D2F0DA000CE178AC;
defparam prom_inst_1.INIT_RAM_1B = 256'hC18D1BF7937DBEF379D9878CC33922C8659DEA3727C8212F9FDE157B73003CFD;
defparam prom_inst_1.INIT_RAM_1C = 256'h2E014948C7133FB6C2640B0ACFD27FB01583D4D9BC37CEB629273F29EC73FF73;
defparam prom_inst_1.INIT_RAM_1D = 256'h07ACDA3BC066C806CC32082062E6294CAFB95FB516DECAB7F7EE726326CE0289;
defparam prom_inst_1.INIT_RAM_1E = 256'h598B35259E9356D9361628AD1B817B13D44D06E044CFB5AE74D3221A93E8A25B;
defparam prom_inst_1.INIT_RAM_1F = 256'hEF4AC6BF9ADDB2EC7B1D4713678ED69D18F330A1424C9A7C461D95D86BB8E2CD;
defparam prom_inst_1.INIT_RAM_20 = 256'h58CB949723619204ACB94D395961A7C83F0532926C5FC08C3DCC4F2F5367A27C;
defparam prom_inst_1.INIT_RAM_21 = 256'h8D7B0D7B609A655864F1E84EA0D03E4D932302699ADCDF94BF5113DB5964CA46;
defparam prom_inst_1.INIT_RAM_22 = 256'hBC3FFC844C8FCC45382CEFEFFB03C4496A3D80FB4ED63DD0B9F10AF66DBE7DCD;
defparam prom_inst_1.INIT_RAM_23 = 256'h36002018784E49EBBC559F5F8715BD8C4FBB27725FB72CDA49B2DB263884F9DE;
defparam prom_inst_1.INIT_RAM_24 = 256'h9B931889B643D9CEF7DC4CAD9C1A89960010296078D2B009860B8A3FB52B1120;
defparam prom_inst_1.INIT_RAM_25 = 256'hAADB18EF17C76DB87233C336F90FA3A123941CA7192B453411E4C79FA57BEA5E;
defparam prom_inst_1.INIT_RAM_26 = 256'h3AC86C114E299F6AD8400F32154122F5CD62E43AECDD40F40023B10C8772F65A;
defparam prom_inst_1.INIT_RAM_27 = 256'h3F6F672910951A71E821C0D6FBE3F99EB227065525C75A3DB67D9FD29CF3599B;
defparam prom_inst_1.INIT_RAM_28 = 256'h5B81064178DDBDC9D4E8085E9D2796A4E316BCE7C90A5C9B211E16118C72CC02;
defparam prom_inst_1.INIT_RAM_29 = 256'hBF634BC2261E3F8B1290A26C5952188190EF0000E163F959C6362DE68E8FEDCB;
defparam prom_inst_1.INIT_RAM_2A = 256'hF54717A184B9FDCB664988EE6E4C51505E1124FD4C82A358AE5194E4BFF23D21;
defparam prom_inst_1.INIT_RAM_2B = 256'hFD821F3C21E84127E5F2F9710F3AF361AE728F638CD7792A78E20AFE68B31B9A;
defparam prom_inst_1.INIT_RAM_2C = 256'h8D27BE0FE974587C8A2D786CDB36CFB7DB3418054E6FC117002C663B3E3C7FF1;
defparam prom_inst_1.INIT_RAM_2D = 256'h272BD0AD3672CFA4300D6E6416E856D612F0A7EB933E2D725DC6244FCED75F3E;
defparam prom_inst_1.INIT_RAM_2E = 256'h264692819200B093000DDF6FE41E00BDB35BE58A3DE1BD6638A8444C085214CD;
defparam prom_inst_1.INIT_RAM_2F = 256'h99B97B6CCC192A67EDD0F07CC5B324C5B60B1FDD6EDBA74E90C5EA39FD661E4D;
defparam prom_inst_1.INIT_RAM_30 = 256'h408DAF19D6DECD7B5E2BC23C217DB24C92D6936CC752FA4EF1C959240B6CCFD9;
defparam prom_inst_1.INIT_RAM_31 = 256'h602F6E5C9E66664982ACC73FAF7E5EF7E4BDBFFA4E53EA6AE13123B04FB2931F;
defparam prom_inst_1.INIT_RAM_32 = 256'h5838BB8428F363067D91E578F420E4111843044A90C1C8F5487B299897607907;
defparam prom_inst_1.INIT_RAM_33 = 256'h8005863B3AE162CAAFC47B89E415886C2122905D88D99983CFA917A8BB8851EE;
defparam prom_inst_1.INIT_RAM_34 = 256'h0AC4388101A05405245386EDDE5696C221C42C08B020F1968EE86CF07B66298D;
defparam prom_inst_1.INIT_RAM_35 = 256'h6ECD6644F46BCAC5F6D2E7B39F6F1039E8020D10384964EE92C9D8048550A142;
defparam prom_inst_1.INIT_RAM_36 = 256'h03C208C5B02818F4CD52A91AEF90D650805F5100BC06EE61A276E7BC9C7B2E09;
defparam prom_inst_1.INIT_RAM_37 = 256'h9092B2B365B95970C99BB36504CE079C2C82AEA2988DA867B0EC3BCAF3556ACE;
defparam prom_inst_1.INIT_RAM_38 = 256'h007AA28BDF45ECC5B7FFBBF064949545454554622CF311852F3724CBE093BC9B;
defparam prom_inst_1.INIT_RAM_39 = 256'hFE56CFD28B080D98F2ACE110333FC1BD9B7681472C15264E6F96B23A87B4D75B;
defparam prom_inst_1.INIT_RAM_3A = 256'h445DB365EFB6B8D562C83231F527CB4952A375AD9F947ECCC9E6F8ED2B133AD1;
defparam prom_inst_1.INIT_RAM_3B = 256'hDB739CE7309EB5F6E77BCE73AAE00C2FA881E33F8F028E638721C346F379934E;
defparam prom_inst_1.INIT_RAM_3C = 256'h5E2213FB8FB76FFBCE5CE77BD373B2E7FFFFDAF7BCE98B2D77FFC6FEEBDCC739;
defparam prom_inst_1.INIT_RAM_3D = 256'hA5B095110A2B7341B03F3354B14402821A5A86211E8A04C9863B66CD06371164;
defparam prom_inst_1.INIT_RAM_3E = 256'h6649B279826D49665BA79977EDDFB981CCF1DDBE7D6332A7349FB6782D1B0022;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFF00000000000000124A3931DFC048CD21C75224E271272893BFB37D920995;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h76030E4F8B41F32380058003C046930A5218350037281206141212B89A9800C2;
defparam prom_inst_2.INIT_RAM_01 = 256'h0026C1A27618CE240547193471259A800A9756AAA8078BF16D2C6D40BE6EEB6D;
defparam prom_inst_2.INIT_RAM_02 = 256'h02228080AA2A7FAAD5003E99B054074800063C890D120187FD7283A4C12372FC;
defparam prom_inst_2.INIT_RAM_03 = 256'hEA18C88046D0357C08317C4DF1F42A956D9CE1F81B7C0A007C451CB00C10A02A;
defparam prom_inst_2.INIT_RAM_04 = 256'h4B29209104A4223E63A04389E67211626471006A9187142976438200115AAA11;
defparam prom_inst_2.INIT_RAM_05 = 256'h618B223468091E438FF6607DCF6259287496181847453CA12A2109680C19C505;
defparam prom_inst_2.INIT_RAM_06 = 256'h0380030024990B61A50CE650E38E1466A109122C5433390A1040AA19CE421111;
defparam prom_inst_2.INIT_RAM_07 = 256'h40B6D9D912ADB7D2AA8555536D068EDB2515C596AAD2B2DF0F5C8CDC54898824;
defparam prom_inst_2.INIT_RAM_08 = 256'h502ACDB7708AA7AF04A16F0C31A03DB64046EA31C00469815C0BAC33EA2A9628;
defparam prom_inst_2.INIT_RAM_09 = 256'h2827E9FC0952C15400024202C251ED6149CA5415E1515F14E45658A8D5A757C1;
defparam prom_inst_2.INIT_RAM_0A = 256'hF8559483485D8D0D369206012032B0A0932824211D2914082C11110B2074A244;
defparam prom_inst_2.INIT_RAM_0B = 256'h7F8F531A337C2F8390C4043A82D520D5B90136D9345A4C1A6486534415BF2F6E;
defparam prom_inst_2.INIT_RAM_0C = 256'hBD64A26AA3EBEB2D74954A72AA1A7C52AD5A0D9740DE37A0E121B302E361C844;
defparam prom_inst_2.INIT_RAM_0D = 256'hA00BB14568028944B7B665262EC80BB5B1114C2DAB88BA422E91493A63569345;
defparam prom_inst_2.INIT_RAM_0E = 256'hFD6165B18A30B4D3A176F6DDE73BBDC867889BB17E2C6218090A2E2EB389A812;
defparam prom_inst_2.INIT_RAM_0F = 256'hC30C2C05850FC322EADC9AE5762C3672CF9A9E7317403683386DF28E7F5CF808;
defparam prom_inst_2.INIT_RAM_10 = 256'h0414997AC33209079B99C304380A11FE937871994CBCA03DE400D848EC6CE824;
defparam prom_inst_2.INIT_RAM_11 = 256'h870184DAEB05D6EBE86F227A1803E4D88E44415E1EA13364682F0C66E04A86D1;
defparam prom_inst_2.INIT_RAM_12 = 256'h3119DE2B20716FE541F69E32D03291E794941A42A63287A348A9C0AEAA520A1E;
defparam prom_inst_2.INIT_RAM_13 = 256'hD184218012482021800514182003CCC00CB2740268015BC0D738D800DC33373F;
defparam prom_inst_2.INIT_RAM_14 = 256'h05081631C773363C9FA2566F8C03E247B88161B06C85214C06C392019C3C7B91;
defparam prom_inst_2.INIT_RAM_15 = 256'hDAB9D6225984128962B33B2EABEC148571DDD7750B2381D9984936092352073B;
defparam prom_inst_2.INIT_RAM_16 = 256'h00000000381EFC000013715B6B976ADFEAE96C00B69F01544111442EE89DD409;
defparam prom_inst_2.INIT_RAM_17 = 256'h0000000000036B11F80406DDDA6FB5006800002064C7E2C600273D8A18800000;
defparam prom_inst_2.INIT_RAM_18 = 256'hAEBFCD2F39FBD642236758A170B84761011045336EE93BE8A98D012DDD3F02D7;
defparam prom_inst_2.INIT_RAM_19 = 256'h80E7BC5E68184570480012032C81260E2C6FF8A81970500A9484544246800346;
defparam prom_inst_2.INIT_RAM_1A = 256'h4205B624100A07014764EBC2832C358E081026620615717C1030430432FFB8C2;
defparam prom_inst_2.INIT_RAM_1B = 256'hFBB39C798DCE309185396B9210001405410C46144145452E9D0BA85E67888261;
defparam prom_inst_2.INIT_RAM_1C = 256'h3C1991B3C1E9D2E179408D56A149002D4243A41CC2C2651C0026326C907E9E33;
defparam prom_inst_2.INIT_RAM_1D = 256'h018103A0809491F0C121B5004888EC6626681D71743F3E80A54A315654BF9B33;
defparam prom_inst_2.INIT_RAM_1E = 256'h0AB00D07860D91F6A18A62D00080168AE20D00A34213846A75C4211AF3EABAC9;
defparam prom_inst_2.INIT_RAM_1F = 256'hF93DAB405801270B70880EC4C7621004042FB04C9A448AAA0928F93F4310E28B;
defparam prom_inst_2.INIT_RAM_20 = 256'hD60652D54700A0DF3648EBD87248E58062448486EF74C756F60014CAC4C1E819;
defparam prom_inst_2.INIT_RAM_21 = 256'hF85ADEB6186B301051A53242E49806053D3504225C5004A33C999950401C5149;
defparam prom_inst_2.INIT_RAM_22 = 256'hA26940722B117609AE10C143A3DDC2C1ABE50022EB68B2016CF37D6C138E155E;
defparam prom_inst_2.INIT_RAM_23 = 256'h0B9B624F61903B2ED502F4B575015AA408AB62A214B26C072D27BA0800412C09;
defparam prom_inst_2.INIT_RAM_24 = 256'h866BDC9C62588AF299EEE7C186CD801B6904034768F00B1119428AC94D8A102D;
defparam prom_inst_2.INIT_RAM_25 = 256'hC75E0EAD9483F651F318B520A9EAB2A70DBBC340F72F470F0C1CBDAD691AE2BC;
defparam prom_inst_2.INIT_RAM_26 = 256'h7D0FCA0146418002808E50BC9966633840C20358F55042F40076E1ECF75EBCD1;
defparam prom_inst_2.INIT_RAM_27 = 256'h475AD40CD025D601296D1C3B2AE00088A4E0D180050030343A0D0A588CA44503;
defparam prom_inst_2.INIT_RAM_28 = 256'h5028842308153D0583936586851481821582EE40618F34EC17C661398E416A3E;
defparam prom_inst_2.INIT_RAM_29 = 256'h2A026A88C180F5141B2B331E36E1800560DA638141595D10060294488E644800;
defparam prom_inst_2.INIT_RAM_2A = 256'h9C29849107CBAC6267817CF9982699CE551D07D6155AD88ECBEDA136951E3DE0;
defparam prom_inst_2.INIT_RAM_2B = 256'h1160100031373C62A27539EFF01C346D61736993D304AEB0281C9251B9A4D0EE;
defparam prom_inst_2.INIT_RAM_2C = 256'hB8476B4A8E59500B21F32E1C24892D97B8B863150E1280B04C6860693D23A32F;
defparam prom_inst_2.INIT_RAM_2D = 256'h692A9E2B9563EA231E1B6EE59818C493F65B26EA3136BA7E784366CD4BB39779;
defparam prom_inst_2.INIT_RAM_2E = 256'h07F680A10C1461FEBF1046862404040C20430969A6005B19B81343370B506703;
defparam prom_inst_2.INIT_RAM_2F = 256'h15087A2228190841A902A06E8522508106109A9F4652D58AB317EA28F10436CD;
defparam prom_inst_2.INIT_RAM_30 = 256'h10F62A59708AB410150A820E001D087C51CE5228C5309B6AA100502C6A620351;
defparam prom_inst_2.INIT_RAM_31 = 256'hB00B4E316A43448D0BA884235AC214AC64294852D5D2E94AB92510582BA13ACA;
defparam prom_inst_2.INIT_RAM_32 = 256'h525DBA35247B42415D04A5583800A008EC02020D80814426C05A550C654220C0;
defparam prom_inst_2.INIT_RAM_33 = 256'h50058F7B32884A4006CA3A81492E930A4125083D308C6C62A93186A7BA2A48EA;
defparam prom_inst_2.INIT_RAM_34 = 256'hAC9742EDD83B7768480554C80A1180D008010A0583A1A9B4028812A05244A2A1;
defparam prom_inst_2.INIT_RAM_35 = 256'h7E8F40F04A52C220641445091B4691454350DF86BF586C6090C8C01B6ADE0BEB;
defparam prom_inst_2.INIT_RAM_36 = 256'h00C5B680214C1483847E3E035902B1C22C48FC5F2851A90638D2FA0737DF3B89;
defparam prom_inst_2.INIT_RAM_37 = 256'hD0AAA1A1410D105881092041408680202EE27CC3D0003C7B21C872C2D4602A2D;
defparam prom_inst_2.INIT_RAM_38 = 256'h3C309080844042BCB555E32CE6D6D7777777776B7D4B5DA6A2B02EEB10A03EA1;
defparam prom_inst_2.INIT_RAM_39 = 256'h53611A9ACA080CC81006B65004A9407385CE4CDCAFC549E14B1ED55A8508850A;
defparam prom_inst_2.INIT_RAM_3A = 256'h0155251D7217D0848C680A35AD32AE66AD5A4103A5A6B4EE8CA34571009BAC2B;
defparam prom_inst_2.INIT_RAM_3B = 256'hDBF39CE7295ED5F6EF7BCEF39CA0DF247E2F5C695452366A244D1244A452A846;
defparam prom_inst_2.INIT_RAM_3C = 256'hC6EAB4A7BACBDC1DFE5CEBFA150DF66BFFFFDC6FDEEA9A8577FEAAFDEDEB7739;
defparam prom_inst_2.INIT_RAM_3D = 256'h958731F575D3E71B39DFBB2837294D2BD418A0768127E9FCF6FEFCD756EB7578;
defparam prom_inst_2.INIT_RAM_3E = 256'h460930B10A1D4546122248C0CB0329088CF5574621C4E3352506B6A4677055A9;
defparam prom_inst_2.INIT_RAM_3F = 256'hFFFF00000000000000040232005D8000443ACB51004021130A8912B109900984;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h1F337CC9F1D55D60400FE6840024A21444883E3323EDC60EE67666C644C41412;
defparam prom_inst_3.INIT_RAM_01 = 256'h09E1C1E9A1DADF6668ABD2639D44A8F4BD6EA006F3FBCFD9F92A6D08DF096935;
defparam prom_inst_3.INIT_RAM_02 = 256'h88280028202A6C6C6C6C53472086C8400040BAB975F400F647A58363C1E22721;
defparam prom_inst_3.INIT_RAM_03 = 256'hC598CDF452D9644A1F7EFCDD89BBEA878E1F01FF35D5B780C0ABDAC1886BC8A2;
defparam prom_inst_3.INIT_RAM_04 = 256'h6DF3C01E00F392915B4045D00375C44174C1B5121D0C0A0E730635CD1A9DD5C3;
defparam prom_inst_3.INIT_RAM_05 = 256'h7AE6EFBB97488118AD97AD45E67EB7FBEE8497166B0A6C389F4CEA576BBB85AD;
defparam prom_inst_3.INIT_RAM_06 = 256'h0100623254D362ED7DCCA67D20820406880765C9AFA2EEDEEFAF17D5BBB66CE6;
defparam prom_inst_3.INIT_RAM_07 = 256'hA0DF7FE54C7BE6E79ACC51991A61335CD91B32A79B95A4044139977CAB6D68A0;
defparam prom_inst_3.INIT_RAM_08 = 256'h88E73A68F818B66BA73D97F4BAEA37DFEEAB930C109DAEA1C4068AA0800CEAC0;
defparam prom_inst_3.INIT_RAM_09 = 256'h464F91A660BD2446729B94BF6CACB672F280182D76A0844BC21BBD1399D57780;
defparam prom_inst_3.INIT_RAM_0A = 256'h54ECBD87A617D09EFF79CE0731F3435D778718F3EB57598CFF0DDDBDF3AD5EA2;
defparam prom_inst_3.INIT_RAM_0B = 256'h4A777D3DBE95EAD2E775438EC6D772AFF3F088F3B915BD7CFD6B65B5C4697DFD;
defparam prom_inst_3.INIT_RAM_0C = 256'h1710DA9E95B2EA5D73AFC0E6C3A4D8ACD71ED7C76E779F71DCC3D714EBA1B3F4;
defparam prom_inst_3.INIT_RAM_0D = 256'hCC4E5EF64006CC05B56887FBA3E46DE95CD87187D9E8EE9A3BA49406B995E89B;
defparam prom_inst_3.INIT_RAM_0E = 256'h83CA27AD44E2F9514FEFC670D6BD5BF5EBFCB7605097F9913A049BBB97D3F37F;
defparam prom_inst_3.INIT_RAM_0F = 256'h7A8C24BE70396DCC738FAC6701705BDB5FDFBCE04EC12BBEBAE08D8E80DD8632;
defparam prom_inst_3.INIT_RAM_10 = 256'h32C4AFE22EB958152F5A260D53202A5C214DBDCF08291021326A2524FD75507A;
defparam prom_inst_3.INIT_RAM_11 = 256'h920B8052EC0F129A101526E22A818CCDAC8748F251800168C4145F29E1385D19;
defparam prom_inst_3.INIT_RAM_12 = 256'h312FB3B820D5C40747DAB88A9D298F22AC198D0E1E8346E5CBA7E04D4B600D04;
defparam prom_inst_3.INIT_RAM_13 = 256'h1E95A2D04400204003820A20E123078007B3710848123AAC182A288344F9AA70;
defparam prom_inst_3.INIT_RAM_14 = 256'hFC848D539E45DF8AA8615ABC9403FB358B20D5215A50B3B72B4E5311B8A0F46E;
defparam prom_inst_3.INIT_RAM_15 = 256'hEBECDADD30161B69B0DD0D7214543A10D42B0A512DA5CAB40A875FA0815FF80A;
defparam prom_inst_3.INIT_RAM_16 = 256'h00000000080A38000028751248044194430C14008012EBEABBBEAFB507432B0F;
defparam prom_inst_3.INIT_RAM_17 = 256'h00000000000449926806039D5F074B803800000030A080C2000E6CC60C800000;
defparam prom_inst_3.INIT_RAM_18 = 256'hCE260C2CA1689395741D55667F4DBE6C2EBFAFFFA7A7AEE9A958246C32824205;
defparam prom_inst_3.INIT_RAM_19 = 256'h80AF5CEC872D98DFD76DE6D524CF057B5E9F2E77D8EE5B50961060621F809674;
defparam prom_inst_3.INIT_RAM_1A = 256'h6D9FDE83EC01CA9C8AFD1A6B0AEDBF5D4921271DE415E37AEB303DCC76CA795D;
defparam prom_inst_3.INIT_RAM_1B = 256'h989F5F7D5EABBF794D7F9AB724DD7DBD9646612DB827ACBCD933519B7BB0C662;
defparam prom_inst_3.INIT_RAM_1C = 256'h3E03D7CBC3E0A56A55FB1573396983DA0A3D6A1B47E0AD267A9CB47F49D6346B;
defparam prom_inst_3.INIT_RAM_1D = 256'h9DF2EADD21B9674A924725C09FB7EECFAE8E4A74B27F7B792E51FD90C1C22FA7;
defparam prom_inst_3.INIT_RAM_1E = 256'h671445DB27DB9ABC2A2AEB7C4ED7EED1B5647D7807FFCD5F79D491A1EB253E49;
defparam prom_inst_3.INIT_RAM_1F = 256'hDE79FE500B3F8E2FB6D62FDFD5FBEBCE5F7E3956EB7CDB4965E04757B25758CB;
defparam prom_inst_3.INIT_RAM_20 = 256'hEE9CDEAAFAFB7BEF42FBC7FB6E7CE9643367ACE055352AFFF3112773BBEBD28B;
defparam prom_inst_3.INIT_RAM_21 = 256'h7AD7355755DD24E8239ECE717F6A5DE3B1FD0E08D66BCF7AFBB817BA7FBD3DEB;
defparam prom_inst_3.INIT_RAM_22 = 256'hFA8843EAE65645BAE411BA552151A152074B8092D6701057D288EAAE57D5C3BC;
defparam prom_inst_3.INIT_RAM_23 = 256'hA040351DC2D5C08087200446FE853C0BDC79DA9DAB328563A8EDBFDCCF470892;
defparam prom_inst_3.INIT_RAM_24 = 256'hDFB6F0D793374D4F53FFC7F74F5E623FA6178DCECA4BBD333FA8E655963FFC94;
defparam prom_inst_3.INIT_RAM_25 = 256'hB6891D103E11FEE7E39CE79A2B82DCD12B79AF9772B22893BABB945FAF2D5FD6;
defparam prom_inst_3.INIT_RAM_26 = 256'hF64A1D4C2491480A7594B81050C0782F1CFBFCD743B7306200AA05F7EBBDA0ED;
defparam prom_inst_3.INIT_RAM_27 = 256'hF3B1DBB7C8F873BA169BD5EA08C83FF29DDE57002B98B012248B8271CBFFFB27;
defparam prom_inst_3.INIT_RAM_28 = 256'h9DC50951BAA36EE923BCBEA6A65CCACF9D2D6C3013DEE5CB7BE22A8CC1F75D0D;
defparam prom_inst_3.INIT_RAM_29 = 256'h3DB48DE376E3E520ADD775B95A6A6A1EDA6DA4044DB44B7FB2D357FE67C45FFE;
defparam prom_inst_3.INIT_RAM_2A = 256'h3AB3E9C3C5852BB56363FBEE5F4F3BFD20395CDFD2BB62BD19DF42FAE5E95696;
defparam prom_inst_3.INIT_RAM_2B = 256'h99FD51F65DA471543C4711550FBD18CA93BBB7B3F4760BFE892AB3BA93C9EBC5;
defparam prom_inst_3.INIT_RAM_2C = 256'hE846AAF2E1D5BF7D73EABEFCFFFFFCD357E73F4886EEC36FC5183C0D1B5537DF;
defparam prom_inst_3.INIT_RAM_2D = 256'hD8E490937D95E7680880CDAB2EC12497215526D1B5F532385A76A75DBFCB55DB;
defparam prom_inst_3.INIT_RAM_2E = 256'hB77AD890FE04DCFFF0676332BD3302639EB99AFEDE14B4BA22FE5452CE54E787;
defparam prom_inst_3.INIT_RAM_2F = 256'hE8EE2EFBDF54FD3D47A97D4CF4F9FA74F2A4A54C557DBB5782D49ECE2AFB83AC;
defparam prom_inst_3.INIT_RAM_30 = 256'h004517DDD2D94D0A4E09F06E04C3F42A79CA531A1F3BC9007D2C4FBCD7BBFB8E;
defparam prom_inst_3.INIT_RAM_31 = 256'h38B2442EC3BC15CECB42F6A739CEF395F5E779CFC9E548B311AE181C31DAB4FB;
defparam prom_inst_3.INIT_RAM_32 = 256'h67D7BD87A6B7AAF18EDC4491B883304C0F41D32DD0766636E898C6A46238B5B0;
defparam prom_inst_3.INIT_RAM_33 = 256'h5007CD5BF7455F9FFBA35D69BC09074AD521142EC904445355B9DA26FD8F4D77;
defparam prom_inst_3.INIT_RAM_34 = 256'h2CFE5FCF9FF332767CD3B59C9B1DCCDA64CC8D9B798051739AE692D892C6A121;
defparam prom_inst_3.INIT_RAM_35 = 256'hB1563799926CE2331FCF85056B9F8C5CBE679C3CB3D4AA1DA9543C1264B1A30B;
defparam prom_inst_3.INIT_RAM_36 = 256'h34DFDE761CB778D7F064323751F1A51F362D26133728374B0E0109210918A48C;
defparam prom_inst_3.INIT_RAM_37 = 256'h407C9B1B369E6D6F6CD81B360F6A4DF0B70515455E9855CD3C4704E20EBD3112;
defparam prom_inst_3.INIT_RAM_38 = 256'h773F36E67E733E7FD8AA77DDF2D26E9F9E93393329419CD052D02ADAA47C5E79;
defparam prom_inst_3.INIT_RAM_39 = 256'hFB278FDA298C2EEB1FF88DD027F261FFDD3F8583E434FFE70EEC8DC88DF39C16;
defparam prom_inst_3.INIT_RAM_3A = 256'hC7EB9EFE5575D0593B9B7841D0BB4F7BF56DB36FC9D71DACA923B650FA8B24F1;
defparam prom_inst_3.INIT_RAM_3B = 256'hDB8C1D07195EE5F60F420EF01CA99986930B6CEFB49E9AEDF3FEF9DA71387971;
defparam prom_inst_3.INIT_RAM_3C = 256'h64345C2E30FDBFFECFC31DC1F6FEF6ADFC19002FDF7771AFF7F06EFBEEF7B555;
defparam prom_inst_3.INIT_RAM_3D = 256'h84CD191A2083612B3153B180118B1048F29D50182002800AD22C24E402221A42;
defparam prom_inst_3.INIT_RAM_3E = 256'h05ED2E25E048BA05ED1F27509D027CE4A24C9D8522E823ABC75A22A1357280C0;
defparam prom_inst_3.INIT_RAM_3F = 256'hFFFF000000000000002DB12F431A819FB808820E93A994EA4077712E868E2172;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'h493AFF1C9BBB9B4B40027CC36A74615C86A0B256B67CD002EA7C7CC444440445;
defparam prom_inst_4.INIT_RAM_01 = 256'hDA51005ED2B2D65641D5ED47B9E700B4C02D987EAC05AA35452622C44020A840;
defparam prom_inst_4.INIT_RAM_02 = 256'h8208888A2A80EC6C6C6C5FFFA0464ECE00C6BF179558013AB820802041A020DB;
defparam prom_inst_4.INIT_RAM_03 = 256'h4F1DD430625D456997FE24653557F160F01FFE008C50A7610CEFC3008439C2A0;
defparam prom_inst_4.INIT_RAM_04 = 256'h8DB3DA83D40183A14B9640D09173C42045012C1B51100B8C664810CB08A588C4;
defparam prom_inst_4.INIT_RAM_05 = 256'hA2E903E7EB0DC011ADB3DF0D8D2376E69A630325200B96B0B628634B7BC40992;
defparam prom_inst_4.INIT_RAM_06 = 256'h6008011016DA6D04D848A45D000017972A89FF71E592564079FDE2C95590783F;
defparam prom_inst_4.INIT_RAM_07 = 256'hC05FEC0CCA1FE960AAC505410E4D0B678A965605BBA40A69CA97C8135AC04422;
defparam prom_inst_4.INIT_RAM_08 = 256'h83DD67FDF9F5B25C2D6B6ACA481827FAA71A0B0018CB4174288C92093DAC948A;
defparam prom_inst_4.INIT_RAM_09 = 256'hC5C2D9F623A928161080108EE344C931350A2845B5A988C69344528E89B021A1;
defparam prom_inst_4.INIT_RAM_0A = 256'hE4C49D81509C448984888062B24F49AC102231D0D12EA818BA199988D144B7AD;
defparam prom_inst_4.INIT_RAM_0B = 256'h012C0040C79DD38AC86EC13E5F18F0F12FA19049F88FD77C17241A85843AEC48;
defparam prom_inst_4.INIT_RAM_0C = 256'hEB10B8E6B47004A28FE8925F08F4375D0E4C1012A268F0222D88000A0DF5246C;
defparam prom_inst_4.INIT_RAM_0D = 256'h4AE58DAA300D44314D179A048E2CEBA48D622A8E1AA3C788D1E12C264187CE86;
defparam prom_inst_4.INIT_RAM_0E = 256'h56BB8380204A6762F1327228A521909845908849258C48F1D68C3511AFD652BC;
defparam prom_inst_4.INIT_RAM_0F = 256'h78D0777BFD10B2218171042FC0B500A0280C530771891E53E63786D55562A895;
defparam prom_inst_4.INIT_RAM_10 = 256'h2C3189369337D14258E5782ED18AAD135A5A1BA0F4ABF09D277428B846C66C18;
defparam prom_inst_4.INIT_RAM_11 = 256'hACCC5F029EBB669179297916DB141336797F5AB94BEEECD7DC89E2C247C5AC56;
defparam prom_inst_4.INIT_RAM_12 = 256'hDE1281582A260159A225911041900E36BDE1BAA1D0F6395634543991B0A5BD8B;
defparam prom_inst_4.INIT_RAM_13 = 256'hB5495000012000608304141451E10A800ABAF507AAB3B62002CFAFA88B1BB82A;
defparam prom_inst_4.INIT_RAM_14 = 256'h80160108059B749002B490096003E6227003305A02B00DA1A0208B11860D5D5D;
defparam prom_inst_4.INIT_RAM_15 = 256'hAEEF98E268430B4D4220201234740EC621D0F4A28012600805829131830563A9;
defparam prom_inst_4.INIT_RAM_16 = 256'h0000000030050600002586259758B469047130012D60510415EAAFCEACA45408;
defparam prom_inst_4.INIT_RAM_17 = 256'h000000000000A2660788243E10B82800440000E00C4628100031913113000000;
defparam prom_inst_4.INIT_RAM_18 = 256'hCCC0F1D2449028A880A82AA2FEBC021C2FEAAFE64AAFEAFDA8197168045088B8;
defparam prom_inst_4.INIT_RAM_19 = 256'h80C3C8B6419ECC5893AD34912CCD27CB169EA866188810C01602220597202444;
defparam prom_inst_4.INIT_RAM_1A = 256'h44DB6DB7A146CC1A7288FCFD390D36EFC1211FFCE98398425B307888408ABC11;
defparam prom_inst_4.INIT_RAM_1B = 256'h997F7EFDFDCB310E411B1C01B4846DB6DB63B32C996E80E8910A42D386496A41;
defparam prom_inst_4.INIT_RAM_1C = 256'h2F112510C9555A484412393BB15B7C401D134F89B30CCC3D458CB237E5558CEB;
defparam prom_inst_4.INIT_RAM_1D = 256'h2E9323ED350D3168DB4EB5E05190FF573E0200F57D181CF8AD5A7A92A1811244;
defparam prom_inst_4.INIT_RAM_1E = 256'h6F34479DA3169899E821E9344786FFE2912FA9FACB21C62F6CD511F3D18DB249;
defparam prom_inst_4.INIT_RAM_1F = 256'hD929BE5019222E6C3FCFE7480D53DF6770F1328816F3C7290042AB20D992C84B;
defparam prom_inst_4.INIT_RAM_20 = 256'h5C8210EAEAE1F90284984B5857708B662A262EB6EC758467359164DB0811298A;
defparam prom_inst_4.INIT_RAM_21 = 256'h02EE2C37601024A058B2486BA1024777836E0E28152BD5FC192FDEB8F885FE30;
defparam prom_inst_4.INIT_RAM_22 = 256'hD42801000023773B6040D951AB0207400EE782A24890FA4818BAD86EE1C7578E;
defparam prom_inst_4.INIT_RAM_23 = 256'h8846B42AF82580100328C0417B875C1FC2DDBA37BEABEDB2850B9E9C40222D44;
defparam prom_inst_4.INIT_RAM_24 = 256'h8A600C8222278E4214844E31800062100F4B89B4080F12B312240669A70D1F90;
defparam prom_inst_4.INIT_RAM_25 = 256'h2D8968AD5A1094BC6110BEB60D50A0259B58621085B80480132C23EC294E4394;
defparam prom_inst_4.INIT_RAM_26 = 256'h3C28D04820A795BAB1983001B35E78E399B39AE0C7EC70E60032DFB9CCF95011;
defparam prom_inst_4.INIT_RAM_27 = 256'h10A1BC810864A8C020A2870F2A9D40EAAD1898A88EB885B66B9E8A71896CF630;
defparam prom_inst_4.INIT_RAM_28 = 256'h56640D839D332326E0830826B7AACDF519A4A9055920408820A66800408A7483;
defparam prom_inst_4.INIT_RAM_29 = 256'h20C60E789174010000622AB91448015B0C00696849C1515600C204586C046B30;
defparam prom_inst_4.INIT_RAM_2A = 256'h82DD6D8820942A05D30440E809F414100010DC84D75EBD2802288724B5013913;
defparam prom_inst_4.INIT_RAM_2B = 256'hF54C59C40966C393AA54BD63F03434E2307A51022074036D85233AD02A7E988B;
defparam prom_inst_4.INIT_RAM_2C = 256'h098528E097E27B124D10AB64DB76D48007276DEC0116D69F87406868413F6B28;
defparam prom_inst_4.INIT_RAM_2D = 256'h11E83C393E604EE855484C778B176497DE5012DB99941A985A6336450A929630;
defparam prom_inst_4.INIT_RAM_2E = 256'h28A4CBB0735B8D4B65D0468D216620FBAF7B0D4144021F842E00102420C04620;
defparam prom_inst_4.INIT_RAM_2F = 256'hB877683FC308E94E89E0AC24313A783130A4402D1102852A886D827731E59409;
defparam prom_inst_4.INIT_RAM_30 = 256'h99058D53FAF5799DDBAC36CD01F578C9146317AAB59E917FADA54727A93FDC13;
defparam prom_inst_4.INIT_RAM_31 = 256'hF0954D12089D460E96C834BBDCF7B9CE67318EE26C6D084AB131A9F814591215;
defparam prom_inst_4.INIT_RAM_32 = 256'h58FA75542203B310A2C6E6AB30915214BD00C53C40328A5E20BB3EEE80197D53;
defparam prom_inst_4.INIT_RAM_33 = 256'h212B9687395462D5522105E1B20509E88FE28002A3698983F7B3C4A875484416;
defparam prom_inst_4.INIT_RAM_34 = 256'hCEE9BD366E4D67B27593EACED57F9EC2C1D824B4F3002110B20E6CF4AA8705BD;
defparam prom_inst_4.INIT_RAM_35 = 256'hC2394768B66DE6C7C5DAFEF1186FE7BEF9BE6CF33461B0BDE3717A491202BCB3;
defparam prom_inst_4.INIT_RAM_36 = 256'hE4DB6DB42C8231F8F67B3D6CE971DE79325F9A64AB1D2FEDB698F5BEEE99370E;
defparam prom_inst_4.INIT_RAM_37 = 256'h8ADFA22245AF9126891E2245588A17DDD844A800963008732CCB25E69B19138E;
defparam prom_inst_4.INIT_RAM_38 = 256'h0721380F3C479CA1BA006B28665658E8E9E67E0010B00024B7372098EADDB8DF;
defparam prom_inst_4.INIT_RAM_39 = 256'h5374CA9AAA94C88B98008183373F959DF936C7632151B67642749AB949747BD4;
defparam prom_inst_4.INIT_RAM_3A = 256'hCC55A7674A56AE1767DDB349FF33EC68B1601E2CCFD73F88A9C3F251D3622E99;
defparam prom_inst_4.INIT_RAM_3B = 256'hDB7E95E739DED5F6E37BCEF381254E2FCD301103E960B26891A4480AD168F97D;
defparam prom_inst_4.INIT_RAM_3C = 256'hB8CAC5A2BEEDDC1DCE5EEDB9E07F76CEFFFDDC6FDFA8AB07F7FEEEF7EF775555;
defparam prom_inst_4.INIT_RAM_3D = 256'h283026E51A68842408A0087186243C800A829601D5842C0700D1401240CC6516;
defparam prom_inst_4.INIT_RAM_3E = 256'h47C93FA0638A7D47D23E2F1D80760060EE89142D20687BA55FA4A6595C011000;
defparam prom_inst_4.INIT_RAM_3F = 256'hFFFF000000000000000FFA33964F89E7BE76BA9FDB5DA9F6ACFBBE3FB9DF49F1;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'hC1DE24BCE20FD7D600007FBA5F68BFFFD3803E5EEA7F940636A4A40484841C57;
defparam prom_inst_5.INIT_RAM_01 = 256'h7071407050EA52F7B9B9BB0EDF1F313C82ADD8DCAFFA0CA1952943A000103838;
defparam prom_inst_5.INIT_RAM_02 = 256'h2A0282820888EC6C6C6C6DF85E121612001EE2099948001A1851317141705051;
defparam prom_inst_5.INIT_RAM_03 = 256'h5D7BC7B9949D929516DAA5541016D800FFE000002429EF232BAEC000ED3FCAA0;
defparam prom_inst_5.INIT_RAM_04 = 256'h7977A4B0259DEE2843CBD6A02273606957A1B780153A02593ADD3EEDDEF7C0E4;
defparam prom_inst_5.INIT_RAM_05 = 256'hC5F22FEF939BA4412923C5812AABE74001602BB67A9FDDFCFF2F7953FFCCA1F9;
defparam prom_inst_5.INIT_RAM_06 = 256'h0008031020410CEAC0DDEEF14554545FA840BF7BF1E2F6CAFBF5C8F19DB3FF3F;
defparam prom_inst_5.INIT_RAM_07 = 256'h208925C8080927F8CCA1004B9FDDD964CFF38EE0CC912B08F8C48ABA5EC00120;
defparam prom_inst_5.INIT_RAM_08 = 256'hF7D53248BCF592D1AF7BE3004501F248BADCFFF760BB08442000C340192F30CE;
defparam prom_inst_5.INIT_RAM_09 = 256'h70745ED7B53C32ABBFF0FFFAF951217D1C232E047DE9E08693F0C08F1F75BFA7;
defparam prom_inst_5.INIT_RAM_0A = 256'h82109B494A0570E1A48F6003BD4BED2F803482FC048B0E4A9ECDDDD2FD123470;
defparam prom_inst_5.INIT_RAM_0B = 256'h808C2AC460C440BF8FD5CDFD0DBA7DFC2B83D8E53EA755DF1BA418C72048270A;
defparam prom_inst_5.INIT_RAM_0C = 256'hE2969DC57D1C00B08F7AF3175D333A564FDF455638B278600580289688E747B4;
defparam prom_inst_5.INIT_RAM_0D = 256'h78D581E384097199080A0A00DA47B69316A1A6DA97B424ED0939AEA57BEF4AEE;
defparam prom_inst_5.INIT_RAM_0E = 256'h4CA4C2529F5F25941B264BAEAD6B55A5C7C6BA49AD0F4D513E9F714145F15E30;
defparam prom_inst_5.INIT_RAM_0F = 256'hACE8240E5F5598EAB85473AA80B02424A82053113183CE6C439EC4B33E66F905;
defparam prom_inst_5.INIT_RAM_10 = 256'h3EAB9B60FFF1FDDABAD3201055EFEC5E7EF63FD0C62B1000AFD67D7DFFD554DB;
defparam prom_inst_5.INIT_RAM_11 = 256'h940D4E82E68940B07A200A0A3BB2088508C7099AC320AA4C850020474B0052FC;
defparam prom_inst_5.INIT_RAM_12 = 256'h11528856EFAE34C10AA4D4E1C3F41A32B7837B308191911A242020E2943A4F7C;
defparam prom_inst_5.INIT_RAM_13 = 256'h3C08456416440000C201062818A1888008BDB9021BDDDABF2E0808BEABCCCAA6;
defparam prom_inst_5.INIT_RAM_14 = 256'hF50D018034AA75444624B50A4803FBE76800981203A009E3240005FEC4035C51;
defparam prom_inst_5.INIT_RAM_15 = 256'hBAABDAC087280BCB082A82056314002209C070080242010287E795DEBD67BC6C;
defparam prom_inst_5.INIT_RAM_16 = 256'h00000000000000000000000000000000000000000000AEAE45FFFAB5041F940F;
defparam prom_inst_5.INIT_RAM_17 = 256'h00000000000000000000001C0F00100000000000002000000000000000000000;
defparam prom_inst_5.INIT_RAM_18 = 256'h66400000600000C8080AAAA07CE6BDFB3AAAAFDDFC0E841347A3315588210040;
defparam prom_inst_5.INIT_RAM_19 = 256'h408B6F9ADBFFFEFFFEA1D7FE007A1BDFE1D7387D12510BFD1E4000903F200104;
defparam prom_inst_5.INIT_RAM_1A = 256'hFF5864EC7FFBF13DAC5FD60DE01FF8AC9039F337BD2442D7FFF82E7860AE9BBE;
defparam prom_inst_5.INIT_RAM_1B = 256'h880378F1F5587FEF4B5AB7E1FFFF6FF8BFFFEB4BFFFAE12FEFDE7D030810BFFD;
defparam prom_inst_5.INIT_RAM_1C = 256'hAC052868C53F52DF8A3E4AAE17C903F030F703AB0C39DE766C7AFCB39F71EAEF;
defparam prom_inst_5.INIT_RAM_1D = 256'h6BBFD5F01F0FFBFEFFFE95A043FEFA556F91C368025A59DF55E3FFEA2364425C;
defparam prom_inst_5.INIT_RAM_1E = 256'h8D7FA1F510E96F01BF900502FA1744F90AC2D607057FA30A61FF172045001000;
defparam prom_inst_5.INIT_RAM_1F = 256'h9140B47FBBFF8460B5AB4C2915895EF889C0D43A72BA75D7F887B6C91CFAC85C;
defparam prom_inst_5.INIT_RAM_20 = 256'h593ABDAEA2AFDF32FC9CFBDECD63DEFAC3164ADB480031A57C9FF8E03FAE1053;
defparam prom_inst_5.INIT_RAM_21 = 256'h91BF987A2BB6697872F3DDFD39F72BC6816B0B9CB57961D9CE5CF7AEEA2EEC62;
defparam prom_inst_5.INIT_RAM_22 = 256'hF1D6BE1111AFDDE15836B6A8F60010775C0E819ED524C9BED38780F425A3E6FD;
defparam prom_inst_5.INIT_RAM_23 = 256'hF3F07B49492D50112ABDCB497FF99D0A327117B9432A85FC40D83DF1FA0AD3F4;
defparam prom_inst_5.INIT_RAM_24 = 256'hA07D22ABCAED2CE3BCAF624A20A3BFD05188F5F4F80EC22ED03903C9E6CFDF89;
defparam prom_inst_5.INIT_RAM_25 = 256'hEFAB288C5F1FF580295D87175245CF03555F1CFEACB015FC57E9684F214E631C;
defparam prom_inst_5.INIT_RAM_26 = 256'hF7E03EF6FEEE2F6CFFE27807C9B3C33232CDFDBD76BD9632006626B14909F48B;
defparam prom_inst_5.INIT_RAM_27 = 256'h87EADBFA39F33EF17693E659D59FFB533E94FAF88BF74F8D1147F5F7BFDF7BFD;
defparam prom_inst_5.INIT_RAM_28 = 256'hCFFF9BD345EAA6FEC8A01350FA0EFEC9EBEDBAAFF7138BBB4C90FF6037BC7E79;
defparam prom_inst_5.INIT_RAM_29 = 256'h95ED1503BD40EBE764DCC443F59F6FE290F570E7B6A2BB2DC1BA8F3E8317D7FC;
defparam prom_inst_5.INIT_RAM_2A = 256'h26964182B2B3F681436E93C06C0922603BB05FB86EA53A11F69246C88A233633;
defparam prom_inst_5.INIT_RAM_2B = 256'hA38FE0FB6618A00FF07BF2C900787053EA76DF2EBD835041D3F02AA2615B1EB9;
defparam prom_inst_5.INIT_RAM_2C = 256'h9B1E791D13BCE9F2C249A965DB76D69AAF21FD163577FECFAC830990D577C232;
defparam prom_inst_5.INIT_RAM_2D = 256'h098757837ADE4C2A30E05DAE56A036D223FC8FE37F7D0131FB6EEFDFEF9F3D0A;
defparam prom_inst_5.INIT_RAM_2E = 256'hACE6FAB4773B0FD36984CF2F6BEE2EFFC7781B937DFABF2867EC1E2CF8CD9D35;
defparam prom_inst_5.INIT_RAM_2F = 256'hBB7F5AFFFBBDE98F138D2E7DBA7CF13A706C8A89001489134C59877F63E9C72D;
defparam prom_inst_5.INIT_RAM_30 = 256'hF51FCF7A5DFDFFFFFF9CBFDD45FA7B9D346337593D9BA5372FBDC727AABFDF33;
defparam prom_inst_5.INIT_RAM_31 = 256'hF0FF5DB37E9DF77F86CB3CF1CC639CC66739CC726C0D2CCAF5398FF93D7F561F;
defparam prom_inst_5.INIT_RAM_32 = 256'h5CFB17AE07ADFB9DEBF5D4FF70F5FE87FDD2E1FDF4BBC3CEF8EBBFCFCC9EF6DF;
defparam prom_inst_5.INIT_RAM_33 = 256'h35E586D155EF72B5426BD7B9FDAFDD09DF55B82B9DE3A3AB7E7FF7BD37AC4F5D;
defparam prom_inst_5.INIT_RAM_34 = 256'h8B690D264FC9553FB7874ACFFF5FDFE3CDF9BCF676070550F21F6CD7F2558B61;
defparam prom_inst_5.INIT_RAM_35 = 256'hC339D76AFE7F7F97E9DAA587BCDF0508AD334C9A3445E2BE8BC57AF9125AE922;
defparam prom_inst_5.INIT_RAM_36 = 256'hBFF864BA6FF9EBD8FC5A2DE4687B31CDD3FDDAECCBD3AA79F5D5F1EEB6D9BB6D;
defparam prom_inst_5.INIT_RAM_37 = 256'hACD26AEBD5873503AB58EBD579AA05D49808098EE7F46EF64F9BF77FDBDA3E5C;
defparam prom_inst_5.INIT_RAM_38 = 256'h8FA1502FB857DDC9BB54C233E414196968654600000400002B3834DDBCDA38D9;
defparam prom_inst_5.INIT_RAM_39 = 256'h525EBA9110602AAB980183816B36D39DDB36ACD32E5BB64E5B2686FC587D2BA4;
defparam prom_inst_5.INIT_RAM_3A = 256'hF6468F667A96870736E6B31BDAAB684952A01B3CEBEFB9CD8B6BBB3BD7136BD7;
defparam prom_inst_5.INIT_RAM_3B = 256'hDB75ADE739DEB5B6E77BCE739DE74E7EED76B3574B47FB7E9DA746EEFDFED57F;
defparam prom_inst_5.INIT_RAM_3C = 256'h010107EBD7AFE3E3EE5EEDB85777B6EF67FCDAB7BFD0D0AFFFFDEEEFEFB6E26D;
defparam prom_inst_5.INIT_RAM_3D = 256'h0200000080040A004400440048008010012000A00040028009000100090080A0;
defparam prom_inst_5.INIT_RAM_3E = 256'h5F5B7BB67BDEED5F52772D42D90B677B88A33517EB50222D57BFEE0204040210;
defparam prom_inst_5.INIT_RAM_3F = 256'hFFFF000000000000000F6AE7DEDB8B76ACB4F3BBDB5DABB38DDB327B49DB8BD8;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h17133C5624CAB161000CEE844AB02046428CAC32B7CCA2CBA1A5A50D0D0D1D71;
defparam prom_inst_6.INIT_RAM_01 = 256'h8F8E018FAF9909C203D688627906C86195716CFE5E0D796D2C04805F7FEFA8E4;
defparam prom_inst_6.INIT_RAM_02 = 256'h00AA802A0282800000007DFFFEDEDFD200D6D201080000040220C000008021AE;
defparam prom_inst_6.INIT_RAM_03 = 256'h0639DCE7F6DA35FFCE683044FCCA41F3000000019FA88CE67E7A7C0198792AA0;
defparam prom_inst_6.INIT_RAM_04 = 256'h49F381990CCF222B5F00591389ED02C046707409A1E706037633D39D398CB599;
defparam prom_inst_6.INIT_RAM_05 = 256'h31CCC3024E79C758E59B24E58422311B2C97BE5EE548349A90BCC00E4E110D84;
defparam prom_inst_6.INIT_RAM_06 = 256'hE4086132596486332CE2510320C31C10888BA4C08F1A0F7C20971F8D63DE21E6;
defparam prom_inst_6.INIT_RAM_07 = 256'h40ADB658E26DB566AA922A334A75077698B7E36EAAC98425C3DEE660294B1886;
defparam prom_inst_6.INIT_RAM_08 = 256'h98C4AB688F7037CEE529062F28FFAB6CDB4C433558DD25C064028A2CF90C662A;
defparam prom_inst_6.INIT_RAM_09 = 256'h41491846616425567397F39363732771BCB0380A3286865A4BA759A64912611A;
defparam prom_inst_6.INIT_RAM_0A = 256'h793209037B0DC38EB2DF7206136320BCDBE040D31D32396B3BEAAAA1D374DCE5;
defparam prom_inst_6.INIT_RAM_0B = 256'h7794B9DE40E45CF84520470C7C1B10C19D9080D1B9B71F1C21B24BE96C2B0667;
defparam prom_inst_6.INIT_RAM_0C = 256'hC61DB8E4127192525B23987BB83A2064B65C61E6E1B45BA6E6BD9BD0BCBC2280;
defparam prom_inst_6.INIT_RAM_0D = 256'hCDE2128E2009C733268409378A44A29AB4718F8B12E0049801241444C3852E82;
defparam prom_inst_6.INIT_RAM_0E = 256'hFCD0CB998F7E25C075EBD8B1B5AD36984DCEAB66BCB578519264938904423301;
defparam prom_inst_6.INIT_RAM_0F = 256'hF1841498E0DE39824588C8934033B336EDB8CB21079F1AC32A3DF7773FAE7FDC;
defparam prom_inst_6.INIT_RAM_10 = 256'hEC10EDBAD339904BB14B7208DB2299004A32D98B0E903029B26D6060664CCE08;
defparam prom_inst_6.INIT_RAM_11 = 256'h7704EE480FD9D4B8DE4C0579B309EC4D8EC76D9CC599316CEF2C250839180B35;
defparam prom_inst_6.INIT_RAM_12 = 256'h24CB1C339B9CF1E41B369EF82D81FD65301905768293F73A6DA0E46EB2E22C3A;
defparam prom_inst_6.INIT_RAM_13 = 256'h25E420E014001800C0850E3031B141000136310E66F15A26DF22816E462AA89F;
defparam prom_inst_6.INIT_RAM_14 = 256'hD08C653DF2ECD74DDFDC53670403E666E4F0513ECA95658C02F39732CF793F62;
defparam prom_inst_6.INIT_RAM_15 = 256'hDBC9BAB41507030B6599D9531124290641996641D9394890CD86070AD5B4A4EE;
defparam prom_inst_6.INIT_RAM_16 = 256'h00000000381FFF00003FFFFFFFFFFFFFFFFFFC01FFFF041011FFFFC050555009;
defparam prom_inst_6.INIT_RAM_17 = 256'h000000000007FFFFFF8E3FE3F0FFEF807C0000E07CDFFFFF003FFFFF1F800000;
defparam prom_inst_6.INIT_RAM_18 = 256'hEEBFFFFF9FFFFE0A820A28A3FD14414D2AAAAFD4500000401100740077DEFFBF;
defparam prom_inst_6.INIT_RAM_19 = 256'h0064D4F181AEDC1DDA7386D0004CC1830345506C5F73197AD41F3E67DF90B7B2;
defparam prom_inst_6.INIT_RAM_1A = 256'h7C35D784654FD77A773DB9BBB76D33925871AF6630B3390F0D30610C5312FA7A;
defparam prom_inst_6.INIT_RAM_1B = 256'hA2AD1B17466DB93824277B3324C4DDB1D36F210C99738F56FD23CF2F65C8AE02;
defparam prom_inst_6.INIT_RAM_1C = 256'h1F1C90F3C5BCDBB99B3A26745CED804D1041BE1884280C07FF6672391CF13E67;
defparam prom_inst_6.INIT_RAM_1D = 256'hF87348E2459DB079D26DCA809F930B45B6E849A5C7212449A6443FC4D3BFD932;
defparam prom_inst_6.INIT_RAM_1E = 256'h161491D34964B92E99D807DBCB8676CE6EC58663C1F59277F6F112BF33FE0800;
defparam prom_inst_6.INIT_RAM_1F = 256'hC69258900F3761B6341355BA47272DEBE45B1EEDDC71C32B092E7F7349957814;
defparam prom_inst_6.INIT_RAM_20 = 256'h226442C9828349D93329652B7418B8E25A4F9852711B933DB27BB3659D66C820;
defparam prom_inst_6.INIT_RAM_21 = 256'h29CE81919E6BB42010A65663E78A910B1ED8087848211B4F34891A61E110A7B9;
defparam prom_inst_6.INIT_RAM_22 = 256'hC7ED4037739677A4E20CFB44204FEF9C879B02EB49BAE75B00F3F32392110B0F;
defparam prom_inst_6.INIT_RAM_23 = 256'h8713F96F4893A3B6D60B74F5888F7EB604CDFADB8C2267B164265ED3C8D9AF72;
defparam prom_inst_6.INIT_RAM_24 = 256'hE5BA59EF67BC9D5ED3B6D964966FA64B38669997EC6819E65BE6806DB76C1CE1;
defparam prom_inst_6.INIT_RAM_25 = 256'hB69D6F3118F2D660B46808BBADFABE844D1C99F2D27E3799DF1A97F4E73FDF77;
defparam prom_inst_6.INIT_RAM_26 = 256'h3BF7F3C0679FEDBA37AF709F3457E10C0047BBC6DB66D27E00AA546C26271875;
defparam prom_inst_6.INIT_RAM_27 = 256'h4D8EDD8D90EEE5D4C02E5A27ACE549EA8CE7C9AA0A38759485224A10813D3673;
defparam prom_inst_6.INIT_RAM_28 = 256'h5CCC8D2A27B12B6642946D89E7384967AD802B1D78EF766C3649A9C8879B7227;
defparam prom_inst_6.INIT_RAM_29 = 256'h6A9E4EBEF1C135CE9BEBBB233739B76F6C5ABFFFFFDD445E83D2B5FB84C44F73;
defparam prom_inst_6.INIT_RAM_2A = 256'h4BB0F3FDFBFBAB3E70AD28D63E365DDE35CC47674746FC84E9659F1654CD59D6;
defparam prom_inst_6.INIT_RAM_2B = 256'hCD3DD0DA90FE1E692C7095E50033185E61A37198779FACF2AF0CE1CC98C86EE7;
defparam prom_inst_6.INIT_RAM_2C = 256'h6704A99A6ECE312B34B2EC9324C93D856C9D27310B9AF278FCE825696A9ADAC5;
defparam prom_inst_6.INIT_RAM_2D = 256'hC2A69FE51C292DAFCF690C6213CF692FC65000EF191608501872306542C256F1;
defparam prom_inst_6.INIT_RAM_2E = 256'h99BD4C5BCFE6796DFFA16248B726264E0460C02DC61E4716161733B3B68776F2;
defparam prom_inst_6.INIT_RAM_2F = 256'h61C4FC310E699838CE08F9ACE1E3C0E1E2B795450023A74F88C186C46887188B;
defparam prom_inst_6.INIT_RAM_30 = 256'h367734C586F12919C969E6430499CD7E498C4B00373ACA6CF8663CB67531319E;
defparam prom_inst_6.INIT_RAM_31 = 256'hF09104E2E9F2048A59F9E3A5295A52B5F4A56B4B58D6A679A1A6B8F872C99071;
defparam prom_inst_6.INIT_RAM_32 = 256'h638D8C630E518273964CE0890893125C3D07973F41E62E3FA0844A3B267275F1;
defparam prom_inst_6.INIT_RAM_33 = 256'h55245B68131C4ECAAD7F2C25CBFBB303476F99767726E6E3B1F3CC938C761CB0;
defparam prom_inst_6.INIT_RAM_34 = 256'h2EB2464C9E9366725C85BB349188481E5CCB8F93CD81F11F92C4B6EE800487A0;
defparam prom_inst_6.INIT_RAM_35 = 256'h12E371B5D9742632672DC0810A070C49D67598AC91D4EA3289C467C6C5CFE20B;
defparam prom_inst_6.INIT_RAM_36 = 256'hB4D5D763398461E2712C972137CF6797255E6D19D670D2431A7059339B792DCD;
defparam prom_inst_6.INIT_RAM_37 = 256'hCD6AB8B972D31C2AE1CAB972C8E2FE7B8267E6414C90941DF97E5C266D345A04;
defparam prom_inst_6.INIT_RAM_38 = 256'h9B2B9364E3723016DCAA9AC4764663B3B3B67B7F7CFBF9FC60D80C41DD685368;
defparam prom_inst_6.INIT_RAM_39 = 256'hAB6BD55C0460088E5AAE8EE1349B3E43450C1DB087FC9921CD1A632843CE8289;
defparam prom_inst_6.INIT_RAM_3A = 256'h3BBB7C91AF88AEDADDA6CB19EA23AD72A54DECF21D1E77C41182CCB0ADD10D7A;
defparam prom_inst_6.INIT_RAM_3B = 256'h3B8B93E8B9C07662E0F8108C1C1DEBEF368D45A9B99E92EB76DDB3D947234323;
defparam prom_inst_6.INIT_RAM_3C = 256'hFEFEFB278C9DFFFFF7E31DC7B788231FE7FFFEFB7FAFFBAFF7FFEE3F8836E76E;
defparam prom_inst_6.INIT_RAM_3D = 256'hFDFFFFFF7FFBF5FFBBFFBBFFB7FF7FEFFEDFFF5FFFBFFD7FF6FFFEFFF6FF7F5F;
defparam prom_inst_6.INIT_RAM_3E = 256'hC12F2853CF3627C13D1194604DC133C998A19D826C89D5A7E364827DFBFBFDEF;
defparam prom_inst_6.INIT_RAM_3F = 256'hFFFF0000000000000039261E7272891A61DBED8924F27899DC4C632906E9BC42;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h328B18492E490203000DA28440801002C24CA434B280B2CB8381810909091923;
defparam prom_inst_7.INIT_RAM_01 = 256'h00000000014909A0065259257906DAC195417AC95E0A29672C4D8000000021AC;
defparam prom_inst_7.INIT_RAM_02 = 256'hAAAA8000AA807FFFFFFFFFFFFFDEDFDE00DFFFDEDFDE00DFFF860E8600078600;
defparam prom_inst_7.INIT_RAM_03 = 256'h0A3088C7F25395FFC90420447DCD2800000000019BA808E6FC3534010C40000A;
defparam prom_inst_7.INIT_RAM_04 = 256'h49E12089044A227BDA005B13AB460060CEF0D00943EF06084477811410529F13;
defparam prom_inst_7.INIT_RAM_05 = 256'h7107E20404784758CC9A64CC8E2251092D90BC7A42456C08A8B588040C3B870D;
defparam prom_inst_7.INIT_RAM_06 = 256'h810001325B2D863364EAD56371860C11808B80891E1A480E41123F0D720240C0;
defparam prom_inst_7.INIT_RAM_07 = 256'h2880029802524A051132AA6E1C32082811B4048D11318C6C8B9EEEE1719B1A84;
defparam prom_inst_7.INIT_RAM_08 = 256'h1B22000187682DA19084066769C380011840483100102488E4668A6CED403353;
defparam prom_inst_7.INIT_RAM_09 = 256'h010C0000601404006017E31981768EC19D94002B230E04DCD9E31B653021053A;
defparam prom_inst_7.INIT_RAM_0A = 256'h833600037981860F36DF1235036629B8C9E060A20C18313195F33331A23068C5;
defparam prom_inst_7.INIT_RAM_0B = 256'h13B99BDEEA508A78452087207899C1E5BF399180E1929A307192C9EA6C63C56F;
defparam prom_inst_7.INIT_RAM_0C = 256'hEC0DA800212096D25C01107B18022170183035FC434AE94EEF1DBBD394DC2280;
defparam prom_inst_7.INIT_RAM_0D = 256'h8002170C28088732648601338040A01B34018D848060A01828063440A6062504;
defparam prom_inst_7.INIT_RAM_0E = 256'hFCF1DB9BAF3E26B0F5EBDAB8B5AD16985D58BB2E99B9780000E0A61804032008;
defparam prom_inst_7.INIT_RAM_0F = 256'h900415B421CE3B826DCDD8B2682397166CB9C922073E0C40281D6B777FA67FDD;
defparam prom_inst_7.INIT_RAM_10 = 256'hE810EDBAD32E800B918956189A201900C932D91B1E811821B029404066444810;
defparam prom_inst_7.INIT_RAM_11 = 256'hF3E4E6C52FD9EAA4EE440F7B151B27988672B49E663B9B2727242548790A1B35;
defparam prom_inst_7.INIT_RAM_12 = 256'h65DB1C63999C71EC59961EF8288154645039073202A1F33A6480A866B6C0383E;
defparam prom_inst_7.INIT_RAM_13 = 256'h20EC69E8040C0070C18102380882E98809B9790CE66124068F628166CE1110BF;
defparam prom_inst_7.INIT_RAM_14 = 256'h500A251DF6EE634DCFDCC72F0E30D8D01050C33E4A9727064673B6224F396B37;
defparam prom_inst_7.INIT_RAM_15 = 256'h35143425350C861B2CBBCB9D8CB04B4E53C92251CB7B519440154692D5AA94C4;
defparam prom_inst_7.INIT_RAM_16 = 256'h2110921148211104104108889042052244844412484950101400001500554186;
defparam prom_inst_7.INIT_RAM_17 = 256'h22222224924892492492493D3F12209084204920854484211042221120822222;
defparam prom_inst_7.INIT_RAM_18 = 256'h888000000000002A880282820040411015555005400104545111441710422489;
defparam prom_inst_7.INIT_RAM_19 = 256'h006434C988B25425491692480024C284830CD02C4F331988700000000E00B510;
defparam prom_inst_7.INIT_RAM_1A = 256'h0A2CB7A0540D536A7735EB96B769219258D0AF6294B1391D14B0530C37347AEA;
defparam prom_inst_7.INIT_RAM_1B = 256'h22251192A328A8A5242568969442B4934921600448134F5010282F6764C88663;
defparam prom_inst_7.INIT_RAM_1C = 256'h189DB1F384BCDBF5992A2650CDB680201052350884240C0FBD6A22619DA1A222;
defparam prom_inst_7.INIT_RAM_1D = 256'hF169592245B490B5C92BDA40CE8B0944B4C041A7C7232485030E254E5AB5CB72;
defparam prom_inst_7.INIT_RAM_1E = 256'h1A22B3535904B526D5C802C9A982292E26C180EBC0D5327356B002D3338E8800;
defparam prom_inst_7.INIT_RAM_1F = 256'hA392C8A0169561D262395490CC2CB5AB848F3EECDC51A282092E7D733B978014;
defparam prom_inst_7.INIT_RAM_20 = 256'h32EE46F44743A0CB332967797288B4804A45B452F90B971CA26A91AC95664860;
defparam prom_inst_7.INIT_RAM_21 = 256'h295A81A3BEE9B410108D5212C698B29D00B504F8409089A724891D115010D3D9;
defparam prom_inst_7.INIT_RAM_22 = 256'hA644003773B732ACA20DEA0C8240000DABBD02E94898E71900937347B2329D0B;
defparam prom_inst_7.INIT_RAM_23 = 256'h0F43A96709B2A234400BE0E1850D6A384EA5E8EA9B226293242E525228F98636;
defparam prom_inst_7.INIT_RAM_24 = 256'hECDA59E567BA9B5E5396C92CB6EF845B796E195784249BC45BC4022D142A1265;
defparam prom_inst_7.INIT_RAM_25 = 256'h590D67B514600241FE288BAD05F038045D1499E2D22C3719CD12939CEF39DEF7;
defparam prom_inst_7.INIT_RAM_26 = 256'h23F3AB80411E689A10A7508F3057A10E1086AB568D52821400AA44682564B876;
defparam prom_inst_7.INIT_RAM_27 = 256'hDA45254D90AED754E0214267840409228464CB82010820818F65402108B51553;
defparam prom_inst_7.INIT_RAM_28 = 256'h5AAA84AB67912156C2946C9955340522A5A48A1829ED22E432D9C5D8275B6AA6;
defparam prom_inst_7.INIT_RAM_29 = 256'h605A0A0EE1C100DE1BABB9662771B0250010DFF9F9441C5A8152B0EB82440D51;
defparam prom_inst_7.INIT_RAM_2A = 256'hCB68B6DDD9620335928D28D236B6DD8801DC0B3741445C84E965B912404D65D5;
defparam prom_inst_7.INIT_RAM_2B = 256'h4534505AB0781E6B8C31A0A70037285161D32898D79F85B3068CD14498A47666;
defparam prom_inst_7.INIT_RAM_2C = 256'h2304A100375E502B34B2C6B36D9B6012698D4730059A7420FCC00441522ACA65;
defparam prom_inst_7.INIT_RAM_2D = 256'h43002FED142B78B3CE650C4411C74DBA564010A2191004701052364442C25049;
defparam prom_inst_7.INIT_RAM_2E = 256'h19BA004287E6516C9FA364DDB740040C0040412CA2064B160C3303B3B28376F2;
defparam prom_inst_7.INIT_RAM_2F = 256'h40887620047B1071C50071C8408140C0A080D5610031224488C1028859021C8B;
defparam prom_inst_7.INIT_RAM_30 = 256'hB6729ADDC6EAA485D569468600188D36CB18CF0A326A40E650C028B67F20238C;
defparam prom_inst_7.INIT_RAM_31 = 256'hA00A88B163204D894B0943AD6B4AD2B5B5A5294B4C88623503EF90D02921126A;
defparam prom_inst_7.INIT_RAM_32 = 256'hF70F4263042146E1490C285A1802A0482805122981456414C046C933222220E1;
defparam prom_inst_7.INIT_RAM_33 = 256'h74044BD41098DC4AA95A12875BEEB703C92D182976A6E6E6A8E10A5382760848;
defparam prom_inst_7.INIT_RAM_34 = 256'h26B646C992B232485D159B324A00003E98530BA10C85F11BA2C8B7AA544D86A0;
defparam prom_inst_7.INIT_RAM_35 = 256'h326721B149D202606231518112448C44565598ACD3C0E022A1D047C2448FE309;
defparam prom_inst_7.INIT_RAM_36 = 256'h12CCB7C3114C41A65164B343128E2592245A6C3BFC70F9229870889199796CDD;
defparam prom_inst_7.INIT_RAM_37 = 256'hC58A90912351080A40889122D042FA6B866006D318A1B04CF13C4A023170EA08;
defparam prom_inst_7.INIT_RAM_38 = 256'hB92A5340C1606096E0AA8A6452C2F696969329000000000060E80A2155886388;
defparam prom_inst_7.INIT_RAM_39 = 256'hA93955491060088CD2AB0EE015897EC74C1C5CF183FD1B23450A2130068EA3A1;
defparam prom_inst_7.INIT_RAM_3A = 256'h3BA955B0A588AE5ADDE6DF19AA22A536AD5FE5F6353CD2A200A24DA52C88872A;
defparam prom_inst_7.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFDE9ED361D4DA9999AA2E932CC9155A351A706;
defparam prom_inst_7.INIT_RAM_3C = 256'h10001B858E1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3D = 256'h0004008002010040000800100100080020002001000800040020200100200004;
defparam prom_inst_7.INIT_RAM_3E = 256'h422D10F28B7646423F20B870C5C3128899E089862D89C4E28062040000004002;
defparam prom_inst_7.INIT_RAM_3F = 256'hFFFF0000000000000030020A7417001C01C9659124B25919CC8C43110F70AC82;

endmodule //VZROM
